magic
tech sky130A
magscale 1 2
timestamp 1730199687
<< nwell >>
rect 1066 97093 318910 97414
rect 1066 96005 318910 96571
rect 1066 94917 318910 95483
rect 1066 93829 318910 94395
rect 1066 92741 318910 93307
rect 1066 91653 318910 92219
rect 1066 90565 318910 91131
rect 1066 89477 318910 90043
rect 1066 88389 318910 88955
rect 1066 87301 318910 87867
rect 1066 86213 318910 86779
rect 1066 85125 318910 85691
rect 1066 84037 318910 84603
rect 1066 82949 318910 83515
rect 1066 81861 318910 82427
rect 1066 80773 318910 81339
rect 1066 79685 318910 80251
rect 1066 78597 318910 79163
rect 1066 77509 318910 78075
rect 1066 76421 318910 76987
rect 1066 75333 318910 75899
rect 1066 74245 318910 74811
rect 1066 73157 318910 73723
rect 1066 72069 318910 72635
rect 1066 70981 318910 71547
rect 1066 69893 318910 70459
rect 1066 68805 318910 69371
rect 1066 67717 318910 68283
rect 1066 66629 318910 67195
rect 1066 65541 318910 66107
rect 1066 64453 318910 65019
rect 1066 63365 318910 63931
rect 1066 62277 318910 62843
rect 1066 61189 318910 61755
rect 1066 60101 318910 60667
rect 1066 59013 318910 59579
rect 1066 57925 318910 58491
rect 1066 56837 318910 57403
rect 1066 55749 318910 56315
rect 1066 54661 318910 55227
rect 1066 53573 318910 54139
rect 1066 52485 318910 53051
rect 1066 51397 318910 51963
rect 1066 50309 318910 50875
rect 1066 49221 318910 49787
rect 1066 48133 318910 48699
rect 1066 47045 318910 47611
rect 1066 45957 318910 46523
rect 1066 44869 318910 45435
rect 1066 43781 318910 44347
rect 1066 42693 318910 43259
rect 1066 41605 318910 42171
rect 1066 40517 318910 41083
rect 1066 39429 318910 39995
rect 1066 38341 318910 38907
rect 1066 37253 318910 37819
rect 1066 36165 318910 36731
rect 1066 35077 318910 35643
rect 1066 33989 318910 34555
rect 1066 32901 318910 33467
rect 1066 31813 318910 32379
rect 1066 30725 318910 31291
rect 1066 29637 318910 30203
rect 1066 28549 318910 29115
rect 1066 27461 318910 28027
rect 1066 26373 318910 26939
rect 1066 25285 318910 25851
rect 1066 24197 318910 24763
rect 1066 23109 318910 23675
rect 1066 22021 318910 22587
rect 1066 20933 318910 21499
rect 1066 19845 318910 20411
rect 1066 18757 318910 19323
rect 1066 17669 318910 18235
rect 1066 16581 318910 17147
rect 1066 15493 318910 16059
rect 1066 14405 318910 14971
rect 1066 13317 318910 13883
rect 1066 12229 318910 12795
rect 1066 11141 318910 11707
rect 1066 10053 318910 10619
rect 1066 8965 318910 9531
rect 1066 7877 318910 8443
rect 1066 6789 318910 7355
rect 1066 5701 318910 6267
rect 1066 4613 318910 5179
rect 1066 3525 318910 4091
rect 1066 2437 318910 3003
<< obsli1 >>
rect 1104 2159 318872 97393
<< obsm1 >>
rect 1104 348 319318 97424
<< metal2 >>
rect 5354 0 5410 800
rect 9770 0 9826 800
rect 14186 0 14242 800
rect 18602 0 18658 800
rect 23018 0 23074 800
rect 27434 0 27490 800
rect 31850 0 31906 800
rect 36266 0 36322 800
rect 40682 0 40738 800
rect 45098 0 45154 800
rect 49514 0 49570 800
rect 53930 0 53986 800
rect 58346 0 58402 800
rect 62762 0 62818 800
rect 67178 0 67234 800
rect 71594 0 71650 800
rect 76010 0 76066 800
rect 80426 0 80482 800
rect 84842 0 84898 800
rect 89258 0 89314 800
rect 93674 0 93730 800
rect 98090 0 98146 800
rect 102506 0 102562 800
rect 106922 0 106978 800
rect 111338 0 111394 800
rect 115754 0 115810 800
rect 120170 0 120226 800
rect 124586 0 124642 800
rect 129002 0 129058 800
rect 133418 0 133474 800
rect 137834 0 137890 800
rect 142250 0 142306 800
rect 146666 0 146722 800
rect 151082 0 151138 800
rect 155498 0 155554 800
rect 159914 0 159970 800
rect 164330 0 164386 800
rect 168746 0 168802 800
rect 173162 0 173218 800
rect 177578 0 177634 800
rect 181994 0 182050 800
rect 186410 0 186466 800
rect 190826 0 190882 800
rect 195242 0 195298 800
rect 199658 0 199714 800
rect 204074 0 204130 800
rect 208490 0 208546 800
rect 212906 0 212962 800
rect 217322 0 217378 800
rect 221738 0 221794 800
rect 226154 0 226210 800
rect 230570 0 230626 800
rect 234986 0 235042 800
rect 239402 0 239458 800
rect 243818 0 243874 800
rect 248234 0 248290 800
rect 252650 0 252706 800
rect 257066 0 257122 800
rect 261482 0 261538 800
rect 265898 0 265954 800
rect 270314 0 270370 800
rect 274730 0 274786 800
rect 279146 0 279202 800
rect 283562 0 283618 800
rect 287978 0 288034 800
rect 292394 0 292450 800
rect 296810 0 296866 800
rect 301226 0 301282 800
rect 305642 0 305698 800
rect 310058 0 310114 800
rect 314474 0 314530 800
<< obsm2 >>
rect 4214 856 319312 98841
rect 4214 342 5298 856
rect 5466 342 9714 856
rect 9882 342 14130 856
rect 14298 342 18546 856
rect 18714 342 22962 856
rect 23130 342 27378 856
rect 27546 342 31794 856
rect 31962 342 36210 856
rect 36378 342 40626 856
rect 40794 342 45042 856
rect 45210 342 49458 856
rect 49626 342 53874 856
rect 54042 342 58290 856
rect 58458 342 62706 856
rect 62874 342 67122 856
rect 67290 342 71538 856
rect 71706 342 75954 856
rect 76122 342 80370 856
rect 80538 342 84786 856
rect 84954 342 89202 856
rect 89370 342 93618 856
rect 93786 342 98034 856
rect 98202 342 102450 856
rect 102618 342 106866 856
rect 107034 342 111282 856
rect 111450 342 115698 856
rect 115866 342 120114 856
rect 120282 342 124530 856
rect 124698 342 128946 856
rect 129114 342 133362 856
rect 133530 342 137778 856
rect 137946 342 142194 856
rect 142362 342 146610 856
rect 146778 342 151026 856
rect 151194 342 155442 856
rect 155610 342 159858 856
rect 160026 342 164274 856
rect 164442 342 168690 856
rect 168858 342 173106 856
rect 173274 342 177522 856
rect 177690 342 181938 856
rect 182106 342 186354 856
rect 186522 342 190770 856
rect 190938 342 195186 856
rect 195354 342 199602 856
rect 199770 342 204018 856
rect 204186 342 208434 856
rect 208602 342 212850 856
rect 213018 342 217266 856
rect 217434 342 221682 856
rect 221850 342 226098 856
rect 226266 342 230514 856
rect 230682 342 234930 856
rect 235098 342 239346 856
rect 239514 342 243762 856
rect 243930 342 248178 856
rect 248346 342 252594 856
rect 252762 342 257010 856
rect 257178 342 261426 856
rect 261594 342 265842 856
rect 266010 342 270258 856
rect 270426 342 274674 856
rect 274842 342 279090 856
rect 279258 342 283506 856
rect 283674 342 287922 856
rect 288090 342 292338 856
rect 292506 342 296754 856
rect 296922 342 301170 856
rect 301338 342 305586 856
rect 305754 342 310002 856
rect 310170 342 314418 856
rect 314586 342 319312 856
<< metal3 >>
rect 319200 98744 320000 98864
rect 319200 96568 320000 96688
rect 319200 94392 320000 94512
rect 319200 92216 320000 92336
rect 319200 90040 320000 90160
rect 319200 87864 320000 87984
rect 319200 85688 320000 85808
rect 319200 83512 320000 83632
rect 319200 81336 320000 81456
rect 319200 79160 320000 79280
rect 319200 76984 320000 77104
rect 319200 74808 320000 74928
rect 319200 72632 320000 72752
rect 319200 70456 320000 70576
rect 319200 68280 320000 68400
rect 319200 66104 320000 66224
rect 319200 63928 320000 64048
rect 319200 61752 320000 61872
rect 319200 59576 320000 59696
rect 319200 57400 320000 57520
rect 319200 55224 320000 55344
rect 319200 53048 320000 53168
rect 319200 50872 320000 50992
rect 319200 48696 320000 48816
rect 319200 46520 320000 46640
rect 319200 44344 320000 44464
rect 319200 42168 320000 42288
rect 319200 39992 320000 40112
rect 319200 37816 320000 37936
rect 319200 35640 320000 35760
rect 319200 33464 320000 33584
rect 319200 31288 320000 31408
rect 319200 29112 320000 29232
rect 319200 26936 320000 27056
rect 319200 24760 320000 24880
rect 319200 22584 320000 22704
rect 319200 20408 320000 20528
rect 319200 18232 320000 18352
rect 319200 16056 320000 16176
rect 319200 13880 320000 14000
rect 319200 11704 320000 11824
rect 319200 9528 320000 9648
rect 319200 7352 320000 7472
rect 319200 5176 320000 5296
rect 319200 3000 320000 3120
rect 319200 824 320000 944
<< obsm3 >>
rect 4210 98664 319120 98837
rect 4210 96768 319227 98664
rect 4210 96488 319120 96768
rect 4210 94592 319227 96488
rect 4210 94312 319120 94592
rect 4210 92416 319227 94312
rect 4210 92136 319120 92416
rect 4210 90240 319227 92136
rect 4210 89960 319120 90240
rect 4210 88064 319227 89960
rect 4210 87784 319120 88064
rect 4210 85888 319227 87784
rect 4210 85608 319120 85888
rect 4210 83712 319227 85608
rect 4210 83432 319120 83712
rect 4210 81536 319227 83432
rect 4210 81256 319120 81536
rect 4210 79360 319227 81256
rect 4210 79080 319120 79360
rect 4210 77184 319227 79080
rect 4210 76904 319120 77184
rect 4210 75008 319227 76904
rect 4210 74728 319120 75008
rect 4210 72832 319227 74728
rect 4210 72552 319120 72832
rect 4210 70656 319227 72552
rect 4210 70376 319120 70656
rect 4210 68480 319227 70376
rect 4210 68200 319120 68480
rect 4210 66304 319227 68200
rect 4210 66024 319120 66304
rect 4210 64128 319227 66024
rect 4210 63848 319120 64128
rect 4210 61952 319227 63848
rect 4210 61672 319120 61952
rect 4210 59776 319227 61672
rect 4210 59496 319120 59776
rect 4210 57600 319227 59496
rect 4210 57320 319120 57600
rect 4210 55424 319227 57320
rect 4210 55144 319120 55424
rect 4210 53248 319227 55144
rect 4210 52968 319120 53248
rect 4210 51072 319227 52968
rect 4210 50792 319120 51072
rect 4210 48896 319227 50792
rect 4210 48616 319120 48896
rect 4210 46720 319227 48616
rect 4210 46440 319120 46720
rect 4210 44544 319227 46440
rect 4210 44264 319120 44544
rect 4210 42368 319227 44264
rect 4210 42088 319120 42368
rect 4210 40192 319227 42088
rect 4210 39912 319120 40192
rect 4210 38016 319227 39912
rect 4210 37736 319120 38016
rect 4210 35840 319227 37736
rect 4210 35560 319120 35840
rect 4210 33664 319227 35560
rect 4210 33384 319120 33664
rect 4210 31488 319227 33384
rect 4210 31208 319120 31488
rect 4210 29312 319227 31208
rect 4210 29032 319120 29312
rect 4210 27136 319227 29032
rect 4210 26856 319120 27136
rect 4210 24960 319227 26856
rect 4210 24680 319120 24960
rect 4210 22784 319227 24680
rect 4210 22504 319120 22784
rect 4210 20608 319227 22504
rect 4210 20328 319120 20608
rect 4210 18432 319227 20328
rect 4210 18152 319120 18432
rect 4210 16256 319227 18152
rect 4210 15976 319120 16256
rect 4210 14080 319227 15976
rect 4210 13800 319120 14080
rect 4210 11904 319227 13800
rect 4210 11624 319120 11904
rect 4210 9728 319227 11624
rect 4210 9448 319120 9728
rect 4210 7552 319227 9448
rect 4210 7272 319120 7552
rect 4210 5376 319227 7272
rect 4210 5096 319120 5376
rect 4210 3200 319227 5096
rect 4210 2920 319120 3200
rect 4210 1024 319227 2920
rect 4210 744 319120 1024
rect 4210 444 319227 744
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
rect 111728 2128 112048 97424
rect 127088 2128 127408 97424
rect 142448 2128 142768 97424
rect 157808 2128 158128 97424
rect 173168 2128 173488 97424
rect 188528 2128 188848 97424
rect 203888 2128 204208 97424
rect 219248 2128 219568 97424
rect 234608 2128 234928 97424
rect 249968 2128 250288 97424
rect 265328 2128 265648 97424
rect 280688 2128 281008 97424
rect 296048 2128 296368 97424
rect 311408 2128 311728 97424
<< obsm4 >>
rect 72923 2048 80928 97205
rect 81408 2048 96288 97205
rect 96768 2048 111648 97205
rect 112128 2048 127008 97205
rect 127488 2048 142368 97205
rect 142848 2048 157728 97205
rect 158208 2048 173088 97205
rect 173568 2048 188448 97205
rect 188928 2048 203808 97205
rect 204288 2048 219168 97205
rect 219648 2048 234528 97205
rect 235008 2048 249888 97205
rect 250368 2048 265248 97205
rect 265728 2048 280608 97205
rect 281088 2048 295968 97205
rect 296448 2048 311328 97205
rect 311808 2048 315869 97205
rect 72923 443 315869 2048
<< labels >>
rlabel metal2 s 168746 0 168802 800 6 a7[0]
port 1 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 a7[10]
port 2 nsew signal output
rlabel metal2 s 217322 0 217378 800 6 a7[11]
port 3 nsew signal output
rlabel metal2 s 221738 0 221794 800 6 a7[12]
port 4 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 a7[13]
port 5 nsew signal output
rlabel metal2 s 230570 0 230626 800 6 a7[14]
port 6 nsew signal output
rlabel metal2 s 234986 0 235042 800 6 a7[15]
port 7 nsew signal output
rlabel metal2 s 239402 0 239458 800 6 a7[16]
port 8 nsew signal output
rlabel metal2 s 243818 0 243874 800 6 a7[17]
port 9 nsew signal output
rlabel metal2 s 248234 0 248290 800 6 a7[18]
port 10 nsew signal output
rlabel metal2 s 252650 0 252706 800 6 a7[19]
port 11 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 a7[1]
port 12 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 a7[20]
port 13 nsew signal output
rlabel metal2 s 261482 0 261538 800 6 a7[21]
port 14 nsew signal output
rlabel metal2 s 265898 0 265954 800 6 a7[22]
port 15 nsew signal output
rlabel metal2 s 270314 0 270370 800 6 a7[23]
port 16 nsew signal output
rlabel metal2 s 274730 0 274786 800 6 a7[24]
port 17 nsew signal output
rlabel metal2 s 279146 0 279202 800 6 a7[25]
port 18 nsew signal output
rlabel metal2 s 283562 0 283618 800 6 a7[26]
port 19 nsew signal output
rlabel metal2 s 287978 0 288034 800 6 a7[27]
port 20 nsew signal output
rlabel metal2 s 292394 0 292450 800 6 a7[28]
port 21 nsew signal output
rlabel metal2 s 296810 0 296866 800 6 a7[29]
port 22 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 a7[2]
port 23 nsew signal output
rlabel metal2 s 301226 0 301282 800 6 a7[30]
port 24 nsew signal output
rlabel metal2 s 305642 0 305698 800 6 a7[31]
port 25 nsew signal output
rlabel metal2 s 181994 0 182050 800 6 a7[3]
port 26 nsew signal output
rlabel metal2 s 186410 0 186466 800 6 a7[4]
port 27 nsew signal output
rlabel metal2 s 190826 0 190882 800 6 a7[5]
port 28 nsew signal output
rlabel metal2 s 195242 0 195298 800 6 a7[6]
port 29 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 a7[7]
port 30 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 a7[8]
port 31 nsew signal output
rlabel metal2 s 208490 0 208546 800 6 a7[9]
port 32 nsew signal output
rlabel metal3 s 319200 824 320000 944 6 csb
port 33 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 gp[0]
port 34 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 gp[10]
port 35 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 gp[11]
port 36 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 gp[12]
port 37 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 gp[13]
port 38 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 gp[14]
port 39 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 gp[15]
port 40 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 gp[16]
port 41 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 gp[17]
port 42 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 gp[18]
port 43 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 gp[19]
port 44 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 gp[1]
port 45 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 gp[20]
port 46 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 gp[21]
port 47 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 gp[22]
port 48 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 gp[23]
port 49 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 gp[24]
port 50 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 gp[25]
port 51 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 gp[26]
port 52 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 gp[27]
port 53 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 gp[28]
port 54 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 gp[29]
port 55 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 gp[2]
port 56 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 gp[30]
port 57 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 gp[31]
port 58 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 gp[3]
port 59 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 gp[4]
port 60 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 gp[5]
port 61 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 gp[6]
port 62 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 gp[7]
port 63 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 gp[8]
port 64 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 gp[9]
port 65 nsew signal output
rlabel metal3 s 319200 81336 320000 81456 6 insMemAddr[0]
port 66 nsew signal output
rlabel metal3 s 319200 83512 320000 83632 6 insMemAddr[1]
port 67 nsew signal output
rlabel metal3 s 319200 85688 320000 85808 6 insMemAddr[2]
port 68 nsew signal output
rlabel metal3 s 319200 87864 320000 87984 6 insMemAddr[3]
port 69 nsew signal output
rlabel metal3 s 319200 90040 320000 90160 6 insMemAddr[4]
port 70 nsew signal output
rlabel metal3 s 319200 92216 320000 92336 6 insMemAddr[5]
port 71 nsew signal output
rlabel metal3 s 319200 94392 320000 94512 6 insMemAddr[6]
port 72 nsew signal output
rlabel metal3 s 319200 96568 320000 96688 6 insMemAddr[7]
port 73 nsew signal output
rlabel metal3 s 319200 98744 320000 98864 6 insMemAddr[8]
port 74 nsew signal output
rlabel metal3 s 319200 11704 320000 11824 6 insMemDataIn[0]
port 75 nsew signal input
rlabel metal3 s 319200 33464 320000 33584 6 insMemDataIn[10]
port 76 nsew signal input
rlabel metal3 s 319200 35640 320000 35760 6 insMemDataIn[11]
port 77 nsew signal input
rlabel metal3 s 319200 37816 320000 37936 6 insMemDataIn[12]
port 78 nsew signal input
rlabel metal3 s 319200 39992 320000 40112 6 insMemDataIn[13]
port 79 nsew signal input
rlabel metal3 s 319200 42168 320000 42288 6 insMemDataIn[14]
port 80 nsew signal input
rlabel metal3 s 319200 44344 320000 44464 6 insMemDataIn[15]
port 81 nsew signal input
rlabel metal3 s 319200 46520 320000 46640 6 insMemDataIn[16]
port 82 nsew signal input
rlabel metal3 s 319200 48696 320000 48816 6 insMemDataIn[17]
port 83 nsew signal input
rlabel metal3 s 319200 50872 320000 50992 6 insMemDataIn[18]
port 84 nsew signal input
rlabel metal3 s 319200 53048 320000 53168 6 insMemDataIn[19]
port 85 nsew signal input
rlabel metal3 s 319200 13880 320000 14000 6 insMemDataIn[1]
port 86 nsew signal input
rlabel metal3 s 319200 55224 320000 55344 6 insMemDataIn[20]
port 87 nsew signal input
rlabel metal3 s 319200 57400 320000 57520 6 insMemDataIn[21]
port 88 nsew signal input
rlabel metal3 s 319200 59576 320000 59696 6 insMemDataIn[22]
port 89 nsew signal input
rlabel metal3 s 319200 61752 320000 61872 6 insMemDataIn[23]
port 90 nsew signal input
rlabel metal3 s 319200 63928 320000 64048 6 insMemDataIn[24]
port 91 nsew signal input
rlabel metal3 s 319200 66104 320000 66224 6 insMemDataIn[25]
port 92 nsew signal input
rlabel metal3 s 319200 68280 320000 68400 6 insMemDataIn[26]
port 93 nsew signal input
rlabel metal3 s 319200 70456 320000 70576 6 insMemDataIn[27]
port 94 nsew signal input
rlabel metal3 s 319200 72632 320000 72752 6 insMemDataIn[28]
port 95 nsew signal input
rlabel metal3 s 319200 74808 320000 74928 6 insMemDataIn[29]
port 96 nsew signal input
rlabel metal3 s 319200 16056 320000 16176 6 insMemDataIn[2]
port 97 nsew signal input
rlabel metal3 s 319200 76984 320000 77104 6 insMemDataIn[30]
port 98 nsew signal input
rlabel metal3 s 319200 79160 320000 79280 6 insMemDataIn[31]
port 99 nsew signal input
rlabel metal3 s 319200 18232 320000 18352 6 insMemDataIn[3]
port 100 nsew signal input
rlabel metal3 s 319200 20408 320000 20528 6 insMemDataIn[4]
port 101 nsew signal input
rlabel metal3 s 319200 22584 320000 22704 6 insMemDataIn[5]
port 102 nsew signal input
rlabel metal3 s 319200 24760 320000 24880 6 insMemDataIn[6]
port 103 nsew signal input
rlabel metal3 s 319200 26936 320000 27056 6 insMemDataIn[7]
port 104 nsew signal input
rlabel metal3 s 319200 29112 320000 29232 6 insMemDataIn[8]
port 105 nsew signal input
rlabel metal3 s 319200 31288 320000 31408 6 insMemDataIn[9]
port 106 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 insMemEn
port 107 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 la_data_in[0]
port 108 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 la_data_in[1]
port 109 nsew signal input
rlabel metal2 s 310058 0 310114 800 6 pc_led
port 110 nsew signal output
rlabel metal2 s 314474 0 314530 800 6 pc_led_oeb
port 111 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 97424 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 97424 6 vssd1
port 113 nsew ground bidirectional
rlabel metal2 s 5354 0 5410 800 6 wb_clk_i
port 114 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wb_rst_i
port 115 nsew signal input
rlabel metal3 s 319200 3000 320000 3120 6 wmask[0]
port 116 nsew signal output
rlabel metal3 s 319200 5176 320000 5296 6 wmask[1]
port 117 nsew signal output
rlabel metal3 s 319200 7352 320000 7472 6 wmask[2]
port 118 nsew signal output
rlabel metal3 s 319200 9528 320000 9648 6 wmask[3]
port 119 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 320000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 69958370
string GDS_FILE /home/jazoolee/uniccass_example/openlane/SLRV/runs/24_10_29_14_34/results/signoff/SLRV.magic.gds
string GDS_START 1654842
<< end >>

