magic
tech sky130A
magscale 1 2
timestamp 1729247982
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 76 558808 349840
<< metal2 >>
rect 3146 0 3202 800
rect 6274 0 6330 800
rect 9402 0 9458 800
rect 12530 0 12586 800
rect 15658 0 15714 800
rect 18786 0 18842 800
rect 21914 0 21970 800
rect 25042 0 25098 800
rect 28170 0 28226 800
rect 31298 0 31354 800
rect 34426 0 34482 800
rect 37554 0 37610 800
rect 40682 0 40738 800
rect 43810 0 43866 800
rect 46938 0 46994 800
rect 50066 0 50122 800
rect 53194 0 53250 800
rect 56322 0 56378 800
rect 59450 0 59506 800
rect 62578 0 62634 800
rect 65706 0 65762 800
rect 68834 0 68890 800
rect 71962 0 72018 800
rect 75090 0 75146 800
rect 78218 0 78274 800
rect 81346 0 81402 800
rect 84474 0 84530 800
rect 87602 0 87658 800
rect 90730 0 90786 800
rect 93858 0 93914 800
rect 96986 0 97042 800
rect 100114 0 100170 800
rect 103242 0 103298 800
rect 106370 0 106426 800
rect 109498 0 109554 800
rect 112626 0 112682 800
rect 115754 0 115810 800
rect 118882 0 118938 800
rect 122010 0 122066 800
rect 125138 0 125194 800
rect 128266 0 128322 800
rect 131394 0 131450 800
rect 134522 0 134578 800
rect 137650 0 137706 800
rect 140778 0 140834 800
rect 143906 0 143962 800
rect 147034 0 147090 800
rect 150162 0 150218 800
rect 153290 0 153346 800
rect 156418 0 156474 800
rect 159546 0 159602 800
rect 162674 0 162730 800
rect 165802 0 165858 800
rect 168930 0 168986 800
rect 172058 0 172114 800
rect 175186 0 175242 800
rect 178314 0 178370 800
rect 181442 0 181498 800
rect 184570 0 184626 800
rect 187698 0 187754 800
rect 190826 0 190882 800
rect 193954 0 194010 800
rect 197082 0 197138 800
rect 200210 0 200266 800
rect 203338 0 203394 800
rect 206466 0 206522 800
rect 209594 0 209650 800
rect 212722 0 212778 800
rect 215850 0 215906 800
rect 218978 0 219034 800
rect 222106 0 222162 800
rect 225234 0 225290 800
rect 228362 0 228418 800
rect 231490 0 231546 800
rect 234618 0 234674 800
rect 237746 0 237802 800
rect 240874 0 240930 800
rect 244002 0 244058 800
rect 247130 0 247186 800
rect 250258 0 250314 800
rect 253386 0 253442 800
rect 256514 0 256570 800
rect 259642 0 259698 800
rect 262770 0 262826 800
rect 265898 0 265954 800
rect 269026 0 269082 800
rect 272154 0 272210 800
rect 275282 0 275338 800
rect 278410 0 278466 800
rect 281538 0 281594 800
rect 284666 0 284722 800
rect 287794 0 287850 800
rect 290922 0 290978 800
rect 294050 0 294106 800
rect 297178 0 297234 800
rect 300306 0 300362 800
rect 303434 0 303490 800
rect 306562 0 306618 800
rect 309690 0 309746 800
rect 312818 0 312874 800
rect 315946 0 316002 800
rect 319074 0 319130 800
rect 322202 0 322258 800
rect 325330 0 325386 800
rect 328458 0 328514 800
rect 331586 0 331642 800
rect 334714 0 334770 800
rect 337842 0 337898 800
rect 340970 0 341026 800
rect 344098 0 344154 800
rect 347226 0 347282 800
rect 350354 0 350410 800
rect 353482 0 353538 800
rect 356610 0 356666 800
rect 359738 0 359794 800
rect 362866 0 362922 800
rect 365994 0 366050 800
rect 369122 0 369178 800
rect 372250 0 372306 800
rect 375378 0 375434 800
rect 378506 0 378562 800
rect 381634 0 381690 800
rect 384762 0 384818 800
rect 387890 0 387946 800
rect 391018 0 391074 800
rect 394146 0 394202 800
rect 397274 0 397330 800
rect 400402 0 400458 800
rect 403530 0 403586 800
rect 406658 0 406714 800
rect 409786 0 409842 800
rect 412914 0 412970 800
rect 416042 0 416098 800
rect 419170 0 419226 800
rect 422298 0 422354 800
rect 425426 0 425482 800
rect 428554 0 428610 800
rect 431682 0 431738 800
rect 434810 0 434866 800
rect 437938 0 437994 800
rect 441066 0 441122 800
rect 444194 0 444250 800
rect 447322 0 447378 800
rect 450450 0 450506 800
rect 453578 0 453634 800
rect 456706 0 456762 800
rect 459834 0 459890 800
rect 462962 0 463018 800
rect 466090 0 466146 800
rect 469218 0 469274 800
rect 472346 0 472402 800
rect 475474 0 475530 800
rect 478602 0 478658 800
rect 481730 0 481786 800
rect 484858 0 484914 800
rect 487986 0 488042 800
rect 491114 0 491170 800
rect 494242 0 494298 800
rect 497370 0 497426 800
rect 500498 0 500554 800
rect 503626 0 503682 800
rect 506754 0 506810 800
rect 509882 0 509938 800
rect 513010 0 513066 800
rect 516138 0 516194 800
rect 519266 0 519322 800
rect 522394 0 522450 800
rect 525522 0 525578 800
rect 528650 0 528706 800
rect 531778 0 531834 800
rect 534906 0 534962 800
rect 538034 0 538090 800
rect 541162 0 541218 800
rect 544290 0 544346 800
rect 547418 0 547474 800
rect 550546 0 550602 800
rect 553674 0 553730 800
rect 556802 0 556858 800
<< obsm2 >>
rect 3148 856 557482 349829
rect 3258 31 6218 856
rect 6386 31 9346 856
rect 9514 31 12474 856
rect 12642 31 15602 856
rect 15770 31 18730 856
rect 18898 31 21858 856
rect 22026 31 24986 856
rect 25154 31 28114 856
rect 28282 31 31242 856
rect 31410 31 34370 856
rect 34538 31 37498 856
rect 37666 31 40626 856
rect 40794 31 43754 856
rect 43922 31 46882 856
rect 47050 31 50010 856
rect 50178 31 53138 856
rect 53306 31 56266 856
rect 56434 31 59394 856
rect 59562 31 62522 856
rect 62690 31 65650 856
rect 65818 31 68778 856
rect 68946 31 71906 856
rect 72074 31 75034 856
rect 75202 31 78162 856
rect 78330 31 81290 856
rect 81458 31 84418 856
rect 84586 31 87546 856
rect 87714 31 90674 856
rect 90842 31 93802 856
rect 93970 31 96930 856
rect 97098 31 100058 856
rect 100226 31 103186 856
rect 103354 31 106314 856
rect 106482 31 109442 856
rect 109610 31 112570 856
rect 112738 31 115698 856
rect 115866 31 118826 856
rect 118994 31 121954 856
rect 122122 31 125082 856
rect 125250 31 128210 856
rect 128378 31 131338 856
rect 131506 31 134466 856
rect 134634 31 137594 856
rect 137762 31 140722 856
rect 140890 31 143850 856
rect 144018 31 146978 856
rect 147146 31 150106 856
rect 150274 31 153234 856
rect 153402 31 156362 856
rect 156530 31 159490 856
rect 159658 31 162618 856
rect 162786 31 165746 856
rect 165914 31 168874 856
rect 169042 31 172002 856
rect 172170 31 175130 856
rect 175298 31 178258 856
rect 178426 31 181386 856
rect 181554 31 184514 856
rect 184682 31 187642 856
rect 187810 31 190770 856
rect 190938 31 193898 856
rect 194066 31 197026 856
rect 197194 31 200154 856
rect 200322 31 203282 856
rect 203450 31 206410 856
rect 206578 31 209538 856
rect 209706 31 212666 856
rect 212834 31 215794 856
rect 215962 31 218922 856
rect 219090 31 222050 856
rect 222218 31 225178 856
rect 225346 31 228306 856
rect 228474 31 231434 856
rect 231602 31 234562 856
rect 234730 31 237690 856
rect 237858 31 240818 856
rect 240986 31 243946 856
rect 244114 31 247074 856
rect 247242 31 250202 856
rect 250370 31 253330 856
rect 253498 31 256458 856
rect 256626 31 259586 856
rect 259754 31 262714 856
rect 262882 31 265842 856
rect 266010 31 268970 856
rect 269138 31 272098 856
rect 272266 31 275226 856
rect 275394 31 278354 856
rect 278522 31 281482 856
rect 281650 31 284610 856
rect 284778 31 287738 856
rect 287906 31 290866 856
rect 291034 31 293994 856
rect 294162 31 297122 856
rect 297290 31 300250 856
rect 300418 31 303378 856
rect 303546 31 306506 856
rect 306674 31 309634 856
rect 309802 31 312762 856
rect 312930 31 315890 856
rect 316058 31 319018 856
rect 319186 31 322146 856
rect 322314 31 325274 856
rect 325442 31 328402 856
rect 328570 31 331530 856
rect 331698 31 334658 856
rect 334826 31 337786 856
rect 337954 31 340914 856
rect 341082 31 344042 856
rect 344210 31 347170 856
rect 347338 31 350298 856
rect 350466 31 353426 856
rect 353594 31 356554 856
rect 356722 31 359682 856
rect 359850 31 362810 856
rect 362978 31 365938 856
rect 366106 31 369066 856
rect 369234 31 372194 856
rect 372362 31 375322 856
rect 375490 31 378450 856
rect 378618 31 381578 856
rect 381746 31 384706 856
rect 384874 31 387834 856
rect 388002 31 390962 856
rect 391130 31 394090 856
rect 394258 31 397218 856
rect 397386 31 400346 856
rect 400514 31 403474 856
rect 403642 31 406602 856
rect 406770 31 409730 856
rect 409898 31 412858 856
rect 413026 31 415986 856
rect 416154 31 419114 856
rect 419282 31 422242 856
rect 422410 31 425370 856
rect 425538 31 428498 856
rect 428666 31 431626 856
rect 431794 31 434754 856
rect 434922 31 437882 856
rect 438050 31 441010 856
rect 441178 31 444138 856
rect 444306 31 447266 856
rect 447434 31 450394 856
rect 450562 31 453522 856
rect 453690 31 456650 856
rect 456818 31 459778 856
rect 459946 31 462906 856
rect 463074 31 466034 856
rect 466202 31 469162 856
rect 469330 31 472290 856
rect 472458 31 475418 856
rect 475586 31 478546 856
rect 478714 31 481674 856
rect 481842 31 484802 856
rect 484970 31 487930 856
rect 488098 31 491058 856
rect 491226 31 494186 856
rect 494354 31 497314 856
rect 497482 31 500442 856
rect 500610 31 503570 856
rect 503738 31 506698 856
rect 506866 31 509826 856
rect 509994 31 512954 856
rect 513122 31 516082 856
rect 516250 31 519210 856
rect 519378 31 522338 856
rect 522506 31 525466 856
rect 525634 31 528594 856
rect 528762 31 531722 856
rect 531890 31 534850 856
rect 535018 31 537978 856
rect 538146 31 541106 856
rect 541274 31 544234 856
rect 544402 31 547362 856
rect 547530 31 550490 856
rect 550658 31 553618 856
rect 553786 31 556746 856
rect 556914 31 557482 856
<< obsm3 >>
rect 4210 35 557486 349825
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 181483 2048 188448 38453
rect 188928 2048 203808 38453
rect 204288 2048 219168 38453
rect 219648 2048 234528 38453
rect 235008 2048 249888 38453
rect 250368 2048 265248 38453
rect 265728 2048 280608 38453
rect 281088 2048 295968 38453
rect 296448 2048 311328 38453
rect 311808 2048 326688 38453
rect 327168 2048 342048 38453
rect 342528 2048 357408 38453
rect 357888 2048 372768 38453
rect 373248 2048 388128 38453
rect 388608 2048 403488 38453
rect 403968 2048 418848 38453
rect 419328 2048 429397 38453
rect 181483 171 429397 2048
<< labels >>
rlabel metal2 s 9402 0 9458 800 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[10]
port 2 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[11]
port 3 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_data_in[12]
port 4 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[13]
port 5 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_data_in[14]
port 6 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[15]
port 7 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[16]
port 8 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[17]
port 9 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_data_in[18]
port 10 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[19]
port 11 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_data_in[1]
port 12 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_data_in[20]
port 13 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[21]
port 14 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[22]
port 15 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[23]
port 16 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_data_in[24]
port 17 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_data_in[25]
port 18 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[26]
port 19 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_data_in[27]
port 20 nsew signal input
rlabel metal2 s 184570 0 184626 800 6 la_data_in[28]
port 21 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_data_in[29]
port 22 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 la_data_in[2]
port 23 nsew signal input
rlabel metal2 s 197082 0 197138 800 6 la_data_in[30]
port 24 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_data_in[31]
port 25 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[32]
port 26 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[33]
port 27 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[34]
port 28 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_data_in[35]
port 29 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_data_in[36]
port 30 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 la_data_in[37]
port 31 nsew signal input
rlabel metal2 s 247130 0 247186 800 6 la_data_in[38]
port 32 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_data_in[39]
port 33 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[3]
port 34 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 la_data_in[40]
port 35 nsew signal input
rlabel metal2 s 265898 0 265954 800 6 la_data_in[41]
port 36 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_data_in[42]
port 37 nsew signal input
rlabel metal2 s 278410 0 278466 800 6 la_data_in[43]
port 38 nsew signal input
rlabel metal2 s 284666 0 284722 800 6 la_data_in[44]
port 39 nsew signal input
rlabel metal2 s 290922 0 290978 800 6 la_data_in[45]
port 40 nsew signal input
rlabel metal2 s 297178 0 297234 800 6 la_data_in[46]
port 41 nsew signal input
rlabel metal2 s 303434 0 303490 800 6 la_data_in[47]
port 42 nsew signal input
rlabel metal2 s 309690 0 309746 800 6 la_data_in[48]
port 43 nsew signal input
rlabel metal2 s 315946 0 316002 800 6 la_data_in[49]
port 44 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[4]
port 45 nsew signal input
rlabel metal2 s 322202 0 322258 800 6 la_data_in[50]
port 46 nsew signal input
rlabel metal2 s 328458 0 328514 800 6 la_data_in[51]
port 47 nsew signal input
rlabel metal2 s 334714 0 334770 800 6 la_data_in[52]
port 48 nsew signal input
rlabel metal2 s 340970 0 341026 800 6 la_data_in[53]
port 49 nsew signal input
rlabel metal2 s 347226 0 347282 800 6 la_data_in[54]
port 50 nsew signal input
rlabel metal2 s 353482 0 353538 800 6 la_data_in[55]
port 51 nsew signal input
rlabel metal2 s 359738 0 359794 800 6 la_data_in[56]
port 52 nsew signal input
rlabel metal2 s 365994 0 366050 800 6 la_data_in[57]
port 53 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 la_data_in[58]
port 54 nsew signal input
rlabel metal2 s 378506 0 378562 800 6 la_data_in[59]
port 55 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_data_in[5]
port 56 nsew signal input
rlabel metal2 s 384762 0 384818 800 6 la_data_in[60]
port 57 nsew signal input
rlabel metal2 s 391018 0 391074 800 6 la_data_in[61]
port 58 nsew signal input
rlabel metal2 s 397274 0 397330 800 6 la_data_in[62]
port 59 nsew signal input
rlabel metal2 s 403530 0 403586 800 6 la_data_in[63]
port 60 nsew signal input
rlabel metal2 s 409786 0 409842 800 6 la_data_in[64]
port 61 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[6]
port 62 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 la_data_in[7]
port 63 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[8]
port 64 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[9]
port 65 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 la_data_out[0]
port 66 nsew signal output
rlabel metal2 s 525522 0 525578 800 6 la_data_out[100]
port 67 nsew signal output
rlabel metal2 s 528650 0 528706 800 6 la_data_out[101]
port 68 nsew signal output
rlabel metal2 s 531778 0 531834 800 6 la_data_out[102]
port 69 nsew signal output
rlabel metal2 s 534906 0 534962 800 6 la_data_out[103]
port 70 nsew signal output
rlabel metal2 s 538034 0 538090 800 6 la_data_out[104]
port 71 nsew signal output
rlabel metal2 s 541162 0 541218 800 6 la_data_out[105]
port 72 nsew signal output
rlabel metal2 s 544290 0 544346 800 6 la_data_out[106]
port 73 nsew signal output
rlabel metal2 s 547418 0 547474 800 6 la_data_out[107]
port 74 nsew signal output
rlabel metal2 s 550546 0 550602 800 6 la_data_out[108]
port 75 nsew signal output
rlabel metal2 s 553674 0 553730 800 6 la_data_out[109]
port 76 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[10]
port 77 nsew signal output
rlabel metal2 s 556802 0 556858 800 6 la_data_out[110]
port 78 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 la_data_out[11]
port 79 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[12]
port 80 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 la_data_out[13]
port 81 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[14]
port 82 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[15]
port 83 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[16]
port 84 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[17]
port 85 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[18]
port 86 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 la_data_out[19]
port 87 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 la_data_out[1]
port 88 nsew signal output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[20]
port 89 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 la_data_out[21]
port 90 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[22]
port 91 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 la_data_out[23]
port 92 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[24]
port 93 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[25]
port 94 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 la_data_out[26]
port 95 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 la_data_out[27]
port 96 nsew signal output
rlabel metal2 s 187698 0 187754 800 6 la_data_out[28]
port 97 nsew signal output
rlabel metal2 s 193954 0 194010 800 6 la_data_out[29]
port 98 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 la_data_out[2]
port 99 nsew signal output
rlabel metal2 s 200210 0 200266 800 6 la_data_out[30]
port 100 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[31]
port 101 nsew signal output
rlabel metal2 s 212722 0 212778 800 6 la_data_out[32]
port 102 nsew signal output
rlabel metal2 s 218978 0 219034 800 6 la_data_out[33]
port 103 nsew signal output
rlabel metal2 s 225234 0 225290 800 6 la_data_out[34]
port 104 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[35]
port 105 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[36]
port 106 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[37]
port 107 nsew signal output
rlabel metal2 s 250258 0 250314 800 6 la_data_out[38]
port 108 nsew signal output
rlabel metal2 s 256514 0 256570 800 6 la_data_out[39]
port 109 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_data_out[3]
port 110 nsew signal output
rlabel metal2 s 262770 0 262826 800 6 la_data_out[40]
port 111 nsew signal output
rlabel metal2 s 269026 0 269082 800 6 la_data_out[41]
port 112 nsew signal output
rlabel metal2 s 275282 0 275338 800 6 la_data_out[42]
port 113 nsew signal output
rlabel metal2 s 281538 0 281594 800 6 la_data_out[43]
port 114 nsew signal output
rlabel metal2 s 287794 0 287850 800 6 la_data_out[44]
port 115 nsew signal output
rlabel metal2 s 294050 0 294106 800 6 la_data_out[45]
port 116 nsew signal output
rlabel metal2 s 300306 0 300362 800 6 la_data_out[46]
port 117 nsew signal output
rlabel metal2 s 306562 0 306618 800 6 la_data_out[47]
port 118 nsew signal output
rlabel metal2 s 312818 0 312874 800 6 la_data_out[48]
port 119 nsew signal output
rlabel metal2 s 319074 0 319130 800 6 la_data_out[49]
port 120 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[4]
port 121 nsew signal output
rlabel metal2 s 325330 0 325386 800 6 la_data_out[50]
port 122 nsew signal output
rlabel metal2 s 331586 0 331642 800 6 la_data_out[51]
port 123 nsew signal output
rlabel metal2 s 337842 0 337898 800 6 la_data_out[52]
port 124 nsew signal output
rlabel metal2 s 344098 0 344154 800 6 la_data_out[53]
port 125 nsew signal output
rlabel metal2 s 350354 0 350410 800 6 la_data_out[54]
port 126 nsew signal output
rlabel metal2 s 356610 0 356666 800 6 la_data_out[55]
port 127 nsew signal output
rlabel metal2 s 362866 0 362922 800 6 la_data_out[56]
port 128 nsew signal output
rlabel metal2 s 369122 0 369178 800 6 la_data_out[57]
port 129 nsew signal output
rlabel metal2 s 375378 0 375434 800 6 la_data_out[58]
port 130 nsew signal output
rlabel metal2 s 381634 0 381690 800 6 la_data_out[59]
port 131 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[5]
port 132 nsew signal output
rlabel metal2 s 387890 0 387946 800 6 la_data_out[60]
port 133 nsew signal output
rlabel metal2 s 394146 0 394202 800 6 la_data_out[61]
port 134 nsew signal output
rlabel metal2 s 400402 0 400458 800 6 la_data_out[62]
port 135 nsew signal output
rlabel metal2 s 406658 0 406714 800 6 la_data_out[63]
port 136 nsew signal output
rlabel metal2 s 412914 0 412970 800 6 la_data_out[64]
port 137 nsew signal output
rlabel metal2 s 416042 0 416098 800 6 la_data_out[65]
port 138 nsew signal output
rlabel metal2 s 419170 0 419226 800 6 la_data_out[66]
port 139 nsew signal output
rlabel metal2 s 422298 0 422354 800 6 la_data_out[67]
port 140 nsew signal output
rlabel metal2 s 425426 0 425482 800 6 la_data_out[68]
port 141 nsew signal output
rlabel metal2 s 428554 0 428610 800 6 la_data_out[69]
port 142 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[6]
port 143 nsew signal output
rlabel metal2 s 431682 0 431738 800 6 la_data_out[70]
port 144 nsew signal output
rlabel metal2 s 434810 0 434866 800 6 la_data_out[71]
port 145 nsew signal output
rlabel metal2 s 437938 0 437994 800 6 la_data_out[72]
port 146 nsew signal output
rlabel metal2 s 441066 0 441122 800 6 la_data_out[73]
port 147 nsew signal output
rlabel metal2 s 444194 0 444250 800 6 la_data_out[74]
port 148 nsew signal output
rlabel metal2 s 447322 0 447378 800 6 la_data_out[75]
port 149 nsew signal output
rlabel metal2 s 450450 0 450506 800 6 la_data_out[76]
port 150 nsew signal output
rlabel metal2 s 453578 0 453634 800 6 la_data_out[77]
port 151 nsew signal output
rlabel metal2 s 456706 0 456762 800 6 la_data_out[78]
port 152 nsew signal output
rlabel metal2 s 459834 0 459890 800 6 la_data_out[79]
port 153 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[7]
port 154 nsew signal output
rlabel metal2 s 462962 0 463018 800 6 la_data_out[80]
port 155 nsew signal output
rlabel metal2 s 466090 0 466146 800 6 la_data_out[81]
port 156 nsew signal output
rlabel metal2 s 469218 0 469274 800 6 la_data_out[82]
port 157 nsew signal output
rlabel metal2 s 472346 0 472402 800 6 la_data_out[83]
port 158 nsew signal output
rlabel metal2 s 475474 0 475530 800 6 la_data_out[84]
port 159 nsew signal output
rlabel metal2 s 478602 0 478658 800 6 la_data_out[85]
port 160 nsew signal output
rlabel metal2 s 481730 0 481786 800 6 la_data_out[86]
port 161 nsew signal output
rlabel metal2 s 484858 0 484914 800 6 la_data_out[87]
port 162 nsew signal output
rlabel metal2 s 487986 0 488042 800 6 la_data_out[88]
port 163 nsew signal output
rlabel metal2 s 491114 0 491170 800 6 la_data_out[89]
port 164 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[8]
port 165 nsew signal output
rlabel metal2 s 494242 0 494298 800 6 la_data_out[90]
port 166 nsew signal output
rlabel metal2 s 497370 0 497426 800 6 la_data_out[91]
port 167 nsew signal output
rlabel metal2 s 500498 0 500554 800 6 la_data_out[92]
port 168 nsew signal output
rlabel metal2 s 503626 0 503682 800 6 la_data_out[93]
port 169 nsew signal output
rlabel metal2 s 506754 0 506810 800 6 la_data_out[94]
port 170 nsew signal output
rlabel metal2 s 509882 0 509938 800 6 la_data_out[95]
port 171 nsew signal output
rlabel metal2 s 513010 0 513066 800 6 la_data_out[96]
port 172 nsew signal output
rlabel metal2 s 516138 0 516194 800 6 la_data_out[97]
port 173 nsew signal output
rlabel metal2 s 519266 0 519322 800 6 la_data_out[98]
port 174 nsew signal output
rlabel metal2 s 522394 0 522450 800 6 la_data_out[99]
port 175 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[9]
port 176 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 178 nsew ground bidirectional
rlabel metal2 s 3146 0 3202 800 6 wb_clk_i
port 179 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wb_rst_i
port 180 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 80197870
string GDS_FILE /home/jazoolee/uniccass_example/openlane/user_proj_example/runs/24_10_18_15_20/results/signoff/user_proj_example.magic.gds
string GDS_START 1267174
<< end >>

