VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SLRV
  CLASS BLOCK ;
  FOREIGN SLRV ;
  ORIGIN 0.000 0.000 ;
  SIZE 1290.000 BY 420.000 ;
  PIN a7[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END a7[0]
  PIN a7[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END a7[10]
  PIN a7[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 877.770 0.000 878.050 4.000 ;
    END
  END a7[11]
  PIN a7[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END a7[12]
  PIN a7[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END a7[13]
  PIN a7[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 931.590 0.000 931.870 4.000 ;
    END
  END a7[14]
  PIN a7[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 4.000 ;
    END
  END a7[15]
  PIN a7[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END a7[16]
  PIN a7[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END a7[17]
  PIN a7[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END a7[18]
  PIN a7[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1021.290 0.000 1021.570 4.000 ;
    END
  END a7[19]
  PIN a7[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END a7[1]
  PIN a7[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1039.230 0.000 1039.510 4.000 ;
    END
  END a7[20]
  PIN a7[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1057.170 0.000 1057.450 4.000 ;
    END
  END a7[21]
  PIN a7[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END a7[22]
  PIN a7[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END a7[23]
  PIN a7[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1110.990 0.000 1111.270 4.000 ;
    END
  END a7[24]
  PIN a7[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END a7[25]
  PIN a7[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1146.870 0.000 1147.150 4.000 ;
    END
  END a7[26]
  PIN a7[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1164.810 0.000 1165.090 4.000 ;
    END
  END a7[27]
  PIN a7[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END a7[28]
  PIN a7[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1200.690 0.000 1200.970 4.000 ;
    END
  END a7[29]
  PIN a7[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END a7[2]
  PIN a7[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1218.630 0.000 1218.910 4.000 ;
    END
  END a7[30]
  PIN a7[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END a7[31]
  PIN a7[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END a7[3]
  PIN a7[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END a7[4]
  PIN a7[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END a7[5]
  PIN a7[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END a7[6]
  PIN a7[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END a7[7]
  PIN a7[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END a7[8]
  PIN a7[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END a7[9]
  PIN csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1286.000 25.880 1290.000 26.480 ;
    END
  END csb
  PIN gp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END gp[0]
  PIN gp[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END gp[10]
  PIN gp[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END gp[11]
  PIN gp[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END gp[12]
  PIN gp[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END gp[13]
  PIN gp[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END gp[14]
  PIN gp[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END gp[15]
  PIN gp[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END gp[16]
  PIN gp[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END gp[17]
  PIN gp[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END gp[18]
  PIN gp[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END gp[19]
  PIN gp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END gp[1]
  PIN gp[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 465.150 0.000 465.430 4.000 ;
    END
  END gp[20]
  PIN gp[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END gp[21]
  PIN gp[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END gp[22]
  PIN gp[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END gp[23]
  PIN gp[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END gp[24]
  PIN gp[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 554.850 0.000 555.130 4.000 ;
    END
  END gp[25]
  PIN gp[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END gp[26]
  PIN gp[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END gp[27]
  PIN gp[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END gp[28]
  PIN gp[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END gp[29]
  PIN gp[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END gp[2]
  PIN gp[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END gp[30]
  PIN gp[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END gp[31]
  PIN gp[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END gp[3]
  PIN gp[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END gp[4]
  PIN gp[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END gp[5]
  PIN gp[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END gp[6]
  PIN gp[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END gp[7]
  PIN gp[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END gp[8]
  PIN gp[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END gp[9]
  PIN insMemAddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 327.800 1290.000 328.400 ;
    END
  END insMemAddr[0]
  PIN insMemAddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 335.960 1290.000 336.560 ;
    END
  END insMemAddr[1]
  PIN insMemAddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 344.120 1290.000 344.720 ;
    END
  END insMemAddr[2]
  PIN insMemAddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 352.280 1290.000 352.880 ;
    END
  END insMemAddr[3]
  PIN insMemAddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 360.440 1290.000 361.040 ;
    END
  END insMemAddr[4]
  PIN insMemAddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 368.600 1290.000 369.200 ;
    END
  END insMemAddr[5]
  PIN insMemAddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 376.760 1290.000 377.360 ;
    END
  END insMemAddr[6]
  PIN insMemAddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 384.920 1290.000 385.520 ;
    END
  END insMemAddr[7]
  PIN insMemAddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 393.080 1290.000 393.680 ;
    END
  END insMemAddr[8]
  PIN insMemDataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 66.680 1290.000 67.280 ;
    END
  END insMemDataIn[0]
  PIN insMemDataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 148.280 1290.000 148.880 ;
    END
  END insMemDataIn[10]
  PIN insMemDataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 156.440 1290.000 157.040 ;
    END
  END insMemDataIn[11]
  PIN insMemDataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 164.600 1290.000 165.200 ;
    END
  END insMemDataIn[12]
  PIN insMemDataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 172.760 1290.000 173.360 ;
    END
  END insMemDataIn[13]
  PIN insMemDataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 180.920 1290.000 181.520 ;
    END
  END insMemDataIn[14]
  PIN insMemDataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 189.080 1290.000 189.680 ;
    END
  END insMemDataIn[15]
  PIN insMemDataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 197.240 1290.000 197.840 ;
    END
  END insMemDataIn[16]
  PIN insMemDataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 205.400 1290.000 206.000 ;
    END
  END insMemDataIn[17]
  PIN insMemDataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 213.560 1290.000 214.160 ;
    END
  END insMemDataIn[18]
  PIN insMemDataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 221.720 1290.000 222.320 ;
    END
  END insMemDataIn[19]
  PIN insMemDataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 74.840 1290.000 75.440 ;
    END
  END insMemDataIn[1]
  PIN insMemDataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 229.880 1290.000 230.480 ;
    END
  END insMemDataIn[20]
  PIN insMemDataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 238.040 1290.000 238.640 ;
    END
  END insMemDataIn[21]
  PIN insMemDataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 246.200 1290.000 246.800 ;
    END
  END insMemDataIn[22]
  PIN insMemDataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 254.360 1290.000 254.960 ;
    END
  END insMemDataIn[23]
  PIN insMemDataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 262.520 1290.000 263.120 ;
    END
  END insMemDataIn[24]
  PIN insMemDataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 270.680 1290.000 271.280 ;
    END
  END insMemDataIn[25]
  PIN insMemDataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 278.840 1290.000 279.440 ;
    END
  END insMemDataIn[26]
  PIN insMemDataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 287.000 1290.000 287.600 ;
    END
  END insMemDataIn[27]
  PIN insMemDataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 295.160 1290.000 295.760 ;
    END
  END insMemDataIn[28]
  PIN insMemDataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 303.320 1290.000 303.920 ;
    END
  END insMemDataIn[29]
  PIN insMemDataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 83.000 1290.000 83.600 ;
    END
  END insMemDataIn[2]
  PIN insMemDataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 311.480 1290.000 312.080 ;
    END
  END insMemDataIn[30]
  PIN insMemDataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 319.640 1290.000 320.240 ;
    END
  END insMemDataIn[31]
  PIN insMemDataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 91.160 1290.000 91.760 ;
    END
  END insMemDataIn[3]
  PIN insMemDataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 99.320 1290.000 99.920 ;
    END
  END insMemDataIn[4]
  PIN insMemDataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 107.480 1290.000 108.080 ;
    END
  END insMemDataIn[5]
  PIN insMemDataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 115.640 1290.000 116.240 ;
    END
  END insMemDataIn[6]
  PIN insMemDataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 123.800 1290.000 124.400 ;
    END
  END insMemDataIn[7]
  PIN insMemDataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 131.960 1290.000 132.560 ;
    END
  END insMemDataIn[8]
  PIN insMemDataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1286.000 140.120 1290.000 140.720 ;
    END
  END insMemDataIn[9]
  PIN insMemEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END insMemEn
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END la_data_in[1]
  PIN pc_led
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1254.510 0.000 1254.790 4.000 ;
    END
  END pc_led
  PIN pc_led_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1272.450 0.000 1272.730 4.000 ;
    END
  END pc_led_oeb
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 408.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 408.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 408.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wb_rst_i
  PIN wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1286.000 34.040 1290.000 34.640 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1286.000 42.200 1290.000 42.800 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1286.000 50.360 1290.000 50.960 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1286.000 58.520 1290.000 59.120 ;
    END
  END wmask[3]
  OBS
      LAYER nwell ;
        RECT 5.330 403.865 1284.510 406.695 ;
        RECT 5.330 398.425 1284.510 401.255 ;
        RECT 5.330 392.985 1284.510 395.815 ;
        RECT 5.330 387.545 1284.510 390.375 ;
        RECT 5.330 382.105 1284.510 384.935 ;
        RECT 5.330 376.665 1284.510 379.495 ;
        RECT 5.330 371.225 1284.510 374.055 ;
        RECT 5.330 365.785 1284.510 368.615 ;
        RECT 5.330 360.345 1284.510 363.175 ;
        RECT 5.330 354.905 1284.510 357.735 ;
        RECT 5.330 349.465 1284.510 352.295 ;
        RECT 5.330 344.025 1284.510 346.855 ;
        RECT 5.330 338.585 1284.510 341.415 ;
        RECT 5.330 333.145 1284.510 335.975 ;
        RECT 5.330 327.705 1284.510 330.535 ;
        RECT 5.330 322.265 1284.510 325.095 ;
        RECT 5.330 316.825 1284.510 319.655 ;
        RECT 5.330 311.385 1284.510 314.215 ;
        RECT 5.330 305.945 1284.510 308.775 ;
        RECT 5.330 300.505 1284.510 303.335 ;
        RECT 5.330 295.065 1284.510 297.895 ;
        RECT 5.330 289.625 1284.510 292.455 ;
        RECT 5.330 284.185 1284.510 287.015 ;
        RECT 5.330 278.745 1284.510 281.575 ;
        RECT 5.330 273.305 1284.510 276.135 ;
        RECT 5.330 267.865 1284.510 270.695 ;
        RECT 5.330 262.425 1284.510 265.255 ;
        RECT 5.330 256.985 1284.510 259.815 ;
        RECT 5.330 251.545 1284.510 254.375 ;
        RECT 5.330 246.105 1284.510 248.935 ;
        RECT 5.330 240.665 1284.510 243.495 ;
        RECT 5.330 235.225 1284.510 238.055 ;
        RECT 5.330 229.785 1284.510 232.615 ;
        RECT 5.330 224.345 1284.510 227.175 ;
        RECT 5.330 218.905 1284.510 221.735 ;
        RECT 5.330 213.465 1284.510 216.295 ;
        RECT 5.330 208.025 1284.510 210.855 ;
        RECT 5.330 202.585 1284.510 205.415 ;
        RECT 5.330 197.145 1284.510 199.975 ;
        RECT 5.330 191.705 1284.510 194.535 ;
        RECT 5.330 186.265 1284.510 189.095 ;
        RECT 5.330 180.825 1284.510 183.655 ;
        RECT 5.330 175.385 1284.510 178.215 ;
        RECT 5.330 169.945 1284.510 172.775 ;
        RECT 5.330 164.505 1284.510 167.335 ;
        RECT 5.330 159.065 1284.510 161.895 ;
        RECT 5.330 153.625 1284.510 156.455 ;
        RECT 5.330 148.185 1284.510 151.015 ;
        RECT 5.330 142.745 1284.510 145.575 ;
        RECT 5.330 137.305 1284.510 140.135 ;
        RECT 5.330 131.865 1284.510 134.695 ;
        RECT 5.330 126.425 1284.510 129.255 ;
        RECT 5.330 120.985 1284.510 123.815 ;
        RECT 5.330 115.545 1284.510 118.375 ;
        RECT 5.330 110.105 1284.510 112.935 ;
        RECT 5.330 104.665 1284.510 107.495 ;
        RECT 5.330 99.225 1284.510 102.055 ;
        RECT 5.330 93.785 1284.510 96.615 ;
        RECT 5.330 88.345 1284.510 91.175 ;
        RECT 5.330 82.905 1284.510 85.735 ;
        RECT 5.330 77.465 1284.510 80.295 ;
        RECT 5.330 72.025 1284.510 74.855 ;
        RECT 5.330 66.585 1284.510 69.415 ;
        RECT 5.330 61.145 1284.510 63.975 ;
        RECT 5.330 55.705 1284.510 58.535 ;
        RECT 5.330 50.265 1284.510 53.095 ;
        RECT 5.330 44.825 1284.510 47.655 ;
        RECT 5.330 39.385 1284.510 42.215 ;
        RECT 5.330 33.945 1284.510 36.775 ;
        RECT 5.330 28.505 1284.510 31.335 ;
        RECT 5.330 23.065 1284.510 25.895 ;
        RECT 5.330 17.625 1284.510 20.455 ;
        RECT 5.330 12.185 1284.510 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1284.320 408.085 ;
      LAYER met1 ;
        RECT 5.520 3.440 1286.090 408.240 ;
      LAYER met2 ;
        RECT 16.660 4.280 1286.060 408.185 ;
        RECT 17.210 2.875 34.310 4.280 ;
        RECT 35.150 2.875 52.250 4.280 ;
        RECT 53.090 2.875 70.190 4.280 ;
        RECT 71.030 2.875 88.130 4.280 ;
        RECT 88.970 2.875 106.070 4.280 ;
        RECT 106.910 2.875 124.010 4.280 ;
        RECT 124.850 2.875 141.950 4.280 ;
        RECT 142.790 2.875 159.890 4.280 ;
        RECT 160.730 2.875 177.830 4.280 ;
        RECT 178.670 2.875 195.770 4.280 ;
        RECT 196.610 2.875 213.710 4.280 ;
        RECT 214.550 2.875 231.650 4.280 ;
        RECT 232.490 2.875 249.590 4.280 ;
        RECT 250.430 2.875 267.530 4.280 ;
        RECT 268.370 2.875 285.470 4.280 ;
        RECT 286.310 2.875 303.410 4.280 ;
        RECT 304.250 2.875 321.350 4.280 ;
        RECT 322.190 2.875 339.290 4.280 ;
        RECT 340.130 2.875 357.230 4.280 ;
        RECT 358.070 2.875 375.170 4.280 ;
        RECT 376.010 2.875 393.110 4.280 ;
        RECT 393.950 2.875 411.050 4.280 ;
        RECT 411.890 2.875 428.990 4.280 ;
        RECT 429.830 2.875 446.930 4.280 ;
        RECT 447.770 2.875 464.870 4.280 ;
        RECT 465.710 2.875 482.810 4.280 ;
        RECT 483.650 2.875 500.750 4.280 ;
        RECT 501.590 2.875 518.690 4.280 ;
        RECT 519.530 2.875 536.630 4.280 ;
        RECT 537.470 2.875 554.570 4.280 ;
        RECT 555.410 2.875 572.510 4.280 ;
        RECT 573.350 2.875 590.450 4.280 ;
        RECT 591.290 2.875 608.390 4.280 ;
        RECT 609.230 2.875 626.330 4.280 ;
        RECT 627.170 2.875 644.270 4.280 ;
        RECT 645.110 2.875 662.210 4.280 ;
        RECT 663.050 2.875 680.150 4.280 ;
        RECT 680.990 2.875 698.090 4.280 ;
        RECT 698.930 2.875 716.030 4.280 ;
        RECT 716.870 2.875 733.970 4.280 ;
        RECT 734.810 2.875 751.910 4.280 ;
        RECT 752.750 2.875 769.850 4.280 ;
        RECT 770.690 2.875 787.790 4.280 ;
        RECT 788.630 2.875 805.730 4.280 ;
        RECT 806.570 2.875 823.670 4.280 ;
        RECT 824.510 2.875 841.610 4.280 ;
        RECT 842.450 2.875 859.550 4.280 ;
        RECT 860.390 2.875 877.490 4.280 ;
        RECT 878.330 2.875 895.430 4.280 ;
        RECT 896.270 2.875 913.370 4.280 ;
        RECT 914.210 2.875 931.310 4.280 ;
        RECT 932.150 2.875 949.250 4.280 ;
        RECT 950.090 2.875 967.190 4.280 ;
        RECT 968.030 2.875 985.130 4.280 ;
        RECT 985.970 2.875 1003.070 4.280 ;
        RECT 1003.910 2.875 1021.010 4.280 ;
        RECT 1021.850 2.875 1038.950 4.280 ;
        RECT 1039.790 2.875 1056.890 4.280 ;
        RECT 1057.730 2.875 1074.830 4.280 ;
        RECT 1075.670 2.875 1092.770 4.280 ;
        RECT 1093.610 2.875 1110.710 4.280 ;
        RECT 1111.550 2.875 1128.650 4.280 ;
        RECT 1129.490 2.875 1146.590 4.280 ;
        RECT 1147.430 2.875 1164.530 4.280 ;
        RECT 1165.370 2.875 1182.470 4.280 ;
        RECT 1183.310 2.875 1200.410 4.280 ;
        RECT 1201.250 2.875 1218.350 4.280 ;
        RECT 1219.190 2.875 1236.290 4.280 ;
        RECT 1237.130 2.875 1254.230 4.280 ;
        RECT 1255.070 2.875 1272.170 4.280 ;
        RECT 1273.010 2.875 1286.060 4.280 ;
      LAYER met3 ;
        RECT 21.050 394.080 1286.000 408.165 ;
        RECT 21.050 392.680 1285.600 394.080 ;
        RECT 21.050 385.920 1286.000 392.680 ;
        RECT 21.050 384.520 1285.600 385.920 ;
        RECT 21.050 377.760 1286.000 384.520 ;
        RECT 21.050 376.360 1285.600 377.760 ;
        RECT 21.050 369.600 1286.000 376.360 ;
        RECT 21.050 368.200 1285.600 369.600 ;
        RECT 21.050 361.440 1286.000 368.200 ;
        RECT 21.050 360.040 1285.600 361.440 ;
        RECT 21.050 353.280 1286.000 360.040 ;
        RECT 21.050 351.880 1285.600 353.280 ;
        RECT 21.050 345.120 1286.000 351.880 ;
        RECT 21.050 343.720 1285.600 345.120 ;
        RECT 21.050 336.960 1286.000 343.720 ;
        RECT 21.050 335.560 1285.600 336.960 ;
        RECT 21.050 328.800 1286.000 335.560 ;
        RECT 21.050 327.400 1285.600 328.800 ;
        RECT 21.050 320.640 1286.000 327.400 ;
        RECT 21.050 319.240 1285.600 320.640 ;
        RECT 21.050 312.480 1286.000 319.240 ;
        RECT 21.050 311.080 1285.600 312.480 ;
        RECT 21.050 304.320 1286.000 311.080 ;
        RECT 21.050 302.920 1285.600 304.320 ;
        RECT 21.050 296.160 1286.000 302.920 ;
        RECT 21.050 294.760 1285.600 296.160 ;
        RECT 21.050 288.000 1286.000 294.760 ;
        RECT 21.050 286.600 1285.600 288.000 ;
        RECT 21.050 279.840 1286.000 286.600 ;
        RECT 21.050 278.440 1285.600 279.840 ;
        RECT 21.050 271.680 1286.000 278.440 ;
        RECT 21.050 270.280 1285.600 271.680 ;
        RECT 21.050 263.520 1286.000 270.280 ;
        RECT 21.050 262.120 1285.600 263.520 ;
        RECT 21.050 255.360 1286.000 262.120 ;
        RECT 21.050 253.960 1285.600 255.360 ;
        RECT 21.050 247.200 1286.000 253.960 ;
        RECT 21.050 245.800 1285.600 247.200 ;
        RECT 21.050 239.040 1286.000 245.800 ;
        RECT 21.050 237.640 1285.600 239.040 ;
        RECT 21.050 230.880 1286.000 237.640 ;
        RECT 21.050 229.480 1285.600 230.880 ;
        RECT 21.050 222.720 1286.000 229.480 ;
        RECT 21.050 221.320 1285.600 222.720 ;
        RECT 21.050 214.560 1286.000 221.320 ;
        RECT 21.050 213.160 1285.600 214.560 ;
        RECT 21.050 206.400 1286.000 213.160 ;
        RECT 21.050 205.000 1285.600 206.400 ;
        RECT 21.050 198.240 1286.000 205.000 ;
        RECT 21.050 196.840 1285.600 198.240 ;
        RECT 21.050 190.080 1286.000 196.840 ;
        RECT 21.050 188.680 1285.600 190.080 ;
        RECT 21.050 181.920 1286.000 188.680 ;
        RECT 21.050 180.520 1285.600 181.920 ;
        RECT 21.050 173.760 1286.000 180.520 ;
        RECT 21.050 172.360 1285.600 173.760 ;
        RECT 21.050 165.600 1286.000 172.360 ;
        RECT 21.050 164.200 1285.600 165.600 ;
        RECT 21.050 157.440 1286.000 164.200 ;
        RECT 21.050 156.040 1285.600 157.440 ;
        RECT 21.050 149.280 1286.000 156.040 ;
        RECT 21.050 147.880 1285.600 149.280 ;
        RECT 21.050 141.120 1286.000 147.880 ;
        RECT 21.050 139.720 1285.600 141.120 ;
        RECT 21.050 132.960 1286.000 139.720 ;
        RECT 21.050 131.560 1285.600 132.960 ;
        RECT 21.050 124.800 1286.000 131.560 ;
        RECT 21.050 123.400 1285.600 124.800 ;
        RECT 21.050 116.640 1286.000 123.400 ;
        RECT 21.050 115.240 1285.600 116.640 ;
        RECT 21.050 108.480 1286.000 115.240 ;
        RECT 21.050 107.080 1285.600 108.480 ;
        RECT 21.050 100.320 1286.000 107.080 ;
        RECT 21.050 98.920 1285.600 100.320 ;
        RECT 21.050 92.160 1286.000 98.920 ;
        RECT 21.050 90.760 1285.600 92.160 ;
        RECT 21.050 84.000 1286.000 90.760 ;
        RECT 21.050 82.600 1285.600 84.000 ;
        RECT 21.050 75.840 1286.000 82.600 ;
        RECT 21.050 74.440 1285.600 75.840 ;
        RECT 21.050 67.680 1286.000 74.440 ;
        RECT 21.050 66.280 1285.600 67.680 ;
        RECT 21.050 59.520 1286.000 66.280 ;
        RECT 21.050 58.120 1285.600 59.520 ;
        RECT 21.050 51.360 1286.000 58.120 ;
        RECT 21.050 49.960 1285.600 51.360 ;
        RECT 21.050 43.200 1286.000 49.960 ;
        RECT 21.050 41.800 1285.600 43.200 ;
        RECT 21.050 35.040 1286.000 41.800 ;
        RECT 21.050 33.640 1285.600 35.040 ;
        RECT 21.050 26.880 1286.000 33.640 ;
        RECT 21.050 25.480 1285.600 26.880 ;
        RECT 21.050 2.895 1286.000 25.480 ;
      LAYER met4 ;
        RECT 132.775 10.240 174.240 390.145 ;
        RECT 176.640 10.240 251.040 390.145 ;
        RECT 253.440 10.240 327.840 390.145 ;
        RECT 330.240 10.240 404.640 390.145 ;
        RECT 407.040 10.240 481.440 390.145 ;
        RECT 483.840 10.240 558.240 390.145 ;
        RECT 560.640 10.240 635.040 390.145 ;
        RECT 637.440 10.240 711.840 390.145 ;
        RECT 714.240 10.240 788.640 390.145 ;
        RECT 791.040 10.240 865.440 390.145 ;
        RECT 867.840 10.240 942.240 390.145 ;
        RECT 944.640 10.240 1019.040 390.145 ;
        RECT 1021.440 10.240 1095.840 390.145 ;
        RECT 1098.240 10.240 1172.640 390.145 ;
        RECT 1175.040 10.240 1249.440 390.145 ;
        RECT 1251.840 10.240 1276.665 390.145 ;
        RECT 132.775 2.895 1276.665 10.240 ;
  END
END SLRV
END LIBRARY

