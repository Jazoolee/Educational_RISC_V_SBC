VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SLRV
  CLASS BLOCK ;
  FOREIGN SLRV ;
  ORIGIN 0.000 0.000 ;
  SIZE 1600.000 BY 500.000 ;
  PIN a7[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END a7[0]
  PIN a7[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1064.530 0.000 1064.810 4.000 ;
    END
  END a7[10]
  PIN a7[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END a7[11]
  PIN a7[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1108.690 0.000 1108.970 4.000 ;
    END
  END a7[12]
  PIN a7[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END a7[13]
  PIN a7[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 0.000 1153.130 4.000 ;
    END
  END a7[14]
  PIN a7[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1174.930 0.000 1175.210 4.000 ;
    END
  END a7[15]
  PIN a7[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1197.010 0.000 1197.290 4.000 ;
    END
  END a7[16]
  PIN a7[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1219.090 0.000 1219.370 4.000 ;
    END
  END a7[17]
  PIN a7[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END a7[18]
  PIN a7[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1263.250 0.000 1263.530 4.000 ;
    END
  END a7[19]
  PIN a7[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END a7[1]
  PIN a7[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1285.330 0.000 1285.610 4.000 ;
    END
  END a7[20]
  PIN a7[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END a7[21]
  PIN a7[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1329.490 0.000 1329.770 4.000 ;
    END
  END a7[22]
  PIN a7[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1351.570 0.000 1351.850 4.000 ;
    END
  END a7[23]
  PIN a7[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1373.650 0.000 1373.930 4.000 ;
    END
  END a7[24]
  PIN a7[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 4.000 ;
    END
  END a7[25]
  PIN a7[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1417.810 0.000 1418.090 4.000 ;
    END
  END a7[26]
  PIN a7[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END a7[27]
  PIN a7[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1461.970 0.000 1462.250 4.000 ;
    END
  END a7[28]
  PIN a7[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1484.050 0.000 1484.330 4.000 ;
    END
  END a7[29]
  PIN a7[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END a7[2]
  PIN a7[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1506.130 0.000 1506.410 4.000 ;
    END
  END a7[30]
  PIN a7[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1528.210 0.000 1528.490 4.000 ;
    END
  END a7[31]
  PIN a7[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 909.970 0.000 910.250 4.000 ;
    END
  END a7[3]
  PIN a7[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END a7[4]
  PIN a7[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 954.130 0.000 954.410 4.000 ;
    END
  END a7[5]
  PIN a7[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END a7[6]
  PIN a7[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END a7[7]
  PIN a7[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END a7[8]
  PIN a7[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1042.450 0.000 1042.730 4.000 ;
    END
  END a7[9]
  PIN csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 4.120 1600.000 4.720 ;
    END
  END csb
  PIN gp[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END gp[0]
  PIN gp[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END gp[10]
  PIN gp[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END gp[11]
  PIN gp[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END gp[12]
  PIN gp[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END gp[13]
  PIN gp[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END gp[14]
  PIN gp[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END gp[15]
  PIN gp[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END gp[16]
  PIN gp[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END gp[17]
  PIN gp[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END gp[18]
  PIN gp[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END gp[19]
  PIN gp[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END gp[1]
  PIN gp[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END gp[20]
  PIN gp[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END gp[21]
  PIN gp[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END gp[22]
  PIN gp[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END gp[23]
  PIN gp[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END gp[24]
  PIN gp[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END gp[25]
  PIN gp[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END gp[26]
  PIN gp[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END gp[27]
  PIN gp[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END gp[28]
  PIN gp[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END gp[29]
  PIN gp[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END gp[2]
  PIN gp[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END gp[30]
  PIN gp[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END gp[31]
  PIN gp[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END gp[3]
  PIN gp[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END gp[4]
  PIN gp[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END gp[5]
  PIN gp[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END gp[6]
  PIN gp[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END gp[7]
  PIN gp[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END gp[8]
  PIN gp[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END gp[9]
  PIN insMemAddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 406.680 1600.000 407.280 ;
    END
  END insMemAddr[0]
  PIN insMemAddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 417.560 1600.000 418.160 ;
    END
  END insMemAddr[1]
  PIN insMemAddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 428.440 1600.000 429.040 ;
    END
  END insMemAddr[2]
  PIN insMemAddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 439.320 1600.000 439.920 ;
    END
  END insMemAddr[3]
  PIN insMemAddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 450.200 1600.000 450.800 ;
    END
  END insMemAddr[4]
  PIN insMemAddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 461.080 1600.000 461.680 ;
    END
  END insMemAddr[5]
  PIN insMemAddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 471.960 1600.000 472.560 ;
    END
  END insMemAddr[6]
  PIN insMemAddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 482.840 1600.000 483.440 ;
    END
  END insMemAddr[7]
  PIN insMemAddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 493.720 1600.000 494.320 ;
    END
  END insMemAddr[8]
  PIN insMemDataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 58.520 1600.000 59.120 ;
    END
  END insMemDataIn[0]
  PIN insMemDataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 167.320 1600.000 167.920 ;
    END
  END insMemDataIn[10]
  PIN insMemDataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 178.200 1600.000 178.800 ;
    END
  END insMemDataIn[11]
  PIN insMemDataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 189.080 1600.000 189.680 ;
    END
  END insMemDataIn[12]
  PIN insMemDataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 199.960 1600.000 200.560 ;
    END
  END insMemDataIn[13]
  PIN insMemDataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 210.840 1600.000 211.440 ;
    END
  END insMemDataIn[14]
  PIN insMemDataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 221.720 1600.000 222.320 ;
    END
  END insMemDataIn[15]
  PIN insMemDataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 232.600 1600.000 233.200 ;
    END
  END insMemDataIn[16]
  PIN insMemDataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 243.480 1600.000 244.080 ;
    END
  END insMemDataIn[17]
  PIN insMemDataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 254.360 1600.000 254.960 ;
    END
  END insMemDataIn[18]
  PIN insMemDataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 265.240 1600.000 265.840 ;
    END
  END insMemDataIn[19]
  PIN insMemDataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 69.400 1600.000 70.000 ;
    END
  END insMemDataIn[1]
  PIN insMemDataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 276.120 1600.000 276.720 ;
    END
  END insMemDataIn[20]
  PIN insMemDataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 287.000 1600.000 287.600 ;
    END
  END insMemDataIn[21]
  PIN insMemDataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 297.880 1600.000 298.480 ;
    END
  END insMemDataIn[22]
  PIN insMemDataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 308.760 1600.000 309.360 ;
    END
  END insMemDataIn[23]
  PIN insMemDataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 319.640 1600.000 320.240 ;
    END
  END insMemDataIn[24]
  PIN insMemDataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 330.520 1600.000 331.120 ;
    END
  END insMemDataIn[25]
  PIN insMemDataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 341.400 1600.000 342.000 ;
    END
  END insMemDataIn[26]
  PIN insMemDataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 352.280 1600.000 352.880 ;
    END
  END insMemDataIn[27]
  PIN insMemDataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 363.160 1600.000 363.760 ;
    END
  END insMemDataIn[28]
  PIN insMemDataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 374.040 1600.000 374.640 ;
    END
  END insMemDataIn[29]
  PIN insMemDataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 80.280 1600.000 80.880 ;
    END
  END insMemDataIn[2]
  PIN insMemDataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 384.920 1600.000 385.520 ;
    END
  END insMemDataIn[30]
  PIN insMemDataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 395.800 1600.000 396.400 ;
    END
  END insMemDataIn[31]
  PIN insMemDataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 91.160 1600.000 91.760 ;
    END
  END insMemDataIn[3]
  PIN insMemDataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 102.040 1600.000 102.640 ;
    END
  END insMemDataIn[4]
  PIN insMemDataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 112.920 1600.000 113.520 ;
    END
  END insMemDataIn[5]
  PIN insMemDataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 123.800 1600.000 124.400 ;
    END
  END insMemDataIn[6]
  PIN insMemDataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 134.680 1600.000 135.280 ;
    END
  END insMemDataIn[7]
  PIN insMemDataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 145.560 1600.000 146.160 ;
    END
  END insMemDataIn[8]
  PIN insMemDataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 1596.000 156.440 1600.000 157.040 ;
    END
  END insMemDataIn[9]
  PIN insMemEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END insMemEn
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END la_data_in[1]
  PIN pc_led
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1550.290 0.000 1550.570 4.000 ;
    END
  END pc_led
  PIN pc_led_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1572.370 0.000 1572.650 4.000 ;
    END
  END pc_led_oeb
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END wb_rst_i
  PIN wmask[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 15.000 1600.000 15.600 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 25.880 1600.000 26.480 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 36.760 1600.000 37.360 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1596.000 47.640 1600.000 48.240 ;
    END
  END wmask[3]
  OBS
      LAYER nwell ;
        RECT 5.330 485.465 1594.550 487.070 ;
        RECT 5.330 480.025 1594.550 482.855 ;
        RECT 5.330 474.585 1594.550 477.415 ;
        RECT 5.330 469.145 1594.550 471.975 ;
        RECT 5.330 463.705 1594.550 466.535 ;
        RECT 5.330 458.265 1594.550 461.095 ;
        RECT 5.330 452.825 1594.550 455.655 ;
        RECT 5.330 447.385 1594.550 450.215 ;
        RECT 5.330 441.945 1594.550 444.775 ;
        RECT 5.330 436.505 1594.550 439.335 ;
        RECT 5.330 431.065 1594.550 433.895 ;
        RECT 5.330 425.625 1594.550 428.455 ;
        RECT 5.330 420.185 1594.550 423.015 ;
        RECT 5.330 414.745 1594.550 417.575 ;
        RECT 5.330 409.305 1594.550 412.135 ;
        RECT 5.330 403.865 1594.550 406.695 ;
        RECT 5.330 398.425 1594.550 401.255 ;
        RECT 5.330 392.985 1594.550 395.815 ;
        RECT 5.330 387.545 1594.550 390.375 ;
        RECT 5.330 382.105 1594.550 384.935 ;
        RECT 5.330 376.665 1594.550 379.495 ;
        RECT 5.330 371.225 1594.550 374.055 ;
        RECT 5.330 365.785 1594.550 368.615 ;
        RECT 5.330 360.345 1594.550 363.175 ;
        RECT 5.330 354.905 1594.550 357.735 ;
        RECT 5.330 349.465 1594.550 352.295 ;
        RECT 5.330 344.025 1594.550 346.855 ;
        RECT 5.330 338.585 1594.550 341.415 ;
        RECT 5.330 333.145 1594.550 335.975 ;
        RECT 5.330 327.705 1594.550 330.535 ;
        RECT 5.330 322.265 1594.550 325.095 ;
        RECT 5.330 316.825 1594.550 319.655 ;
        RECT 5.330 311.385 1594.550 314.215 ;
        RECT 5.330 305.945 1594.550 308.775 ;
        RECT 5.330 300.505 1594.550 303.335 ;
        RECT 5.330 295.065 1594.550 297.895 ;
        RECT 5.330 289.625 1594.550 292.455 ;
        RECT 5.330 284.185 1594.550 287.015 ;
        RECT 5.330 278.745 1594.550 281.575 ;
        RECT 5.330 273.305 1594.550 276.135 ;
        RECT 5.330 267.865 1594.550 270.695 ;
        RECT 5.330 262.425 1594.550 265.255 ;
        RECT 5.330 256.985 1594.550 259.815 ;
        RECT 5.330 251.545 1594.550 254.375 ;
        RECT 5.330 246.105 1594.550 248.935 ;
        RECT 5.330 240.665 1594.550 243.495 ;
        RECT 5.330 235.225 1594.550 238.055 ;
        RECT 5.330 229.785 1594.550 232.615 ;
        RECT 5.330 224.345 1594.550 227.175 ;
        RECT 5.330 218.905 1594.550 221.735 ;
        RECT 5.330 213.465 1594.550 216.295 ;
        RECT 5.330 208.025 1594.550 210.855 ;
        RECT 5.330 202.585 1594.550 205.415 ;
        RECT 5.330 197.145 1594.550 199.975 ;
        RECT 5.330 191.705 1594.550 194.535 ;
        RECT 5.330 186.265 1594.550 189.095 ;
        RECT 5.330 180.825 1594.550 183.655 ;
        RECT 5.330 175.385 1594.550 178.215 ;
        RECT 5.330 169.945 1594.550 172.775 ;
        RECT 5.330 164.505 1594.550 167.335 ;
        RECT 5.330 159.065 1594.550 161.895 ;
        RECT 5.330 153.625 1594.550 156.455 ;
        RECT 5.330 148.185 1594.550 151.015 ;
        RECT 5.330 142.745 1594.550 145.575 ;
        RECT 5.330 137.305 1594.550 140.135 ;
        RECT 5.330 131.865 1594.550 134.695 ;
        RECT 5.330 126.425 1594.550 129.255 ;
        RECT 5.330 120.985 1594.550 123.815 ;
        RECT 5.330 115.545 1594.550 118.375 ;
        RECT 5.330 110.105 1594.550 112.935 ;
        RECT 5.330 104.665 1594.550 107.495 ;
        RECT 5.330 99.225 1594.550 102.055 ;
        RECT 5.330 93.785 1594.550 96.615 ;
        RECT 5.330 88.345 1594.550 91.175 ;
        RECT 5.330 82.905 1594.550 85.735 ;
        RECT 5.330 77.465 1594.550 80.295 ;
        RECT 5.330 72.025 1594.550 74.855 ;
        RECT 5.330 66.585 1594.550 69.415 ;
        RECT 5.330 61.145 1594.550 63.975 ;
        RECT 5.330 55.705 1594.550 58.535 ;
        RECT 5.330 50.265 1594.550 53.095 ;
        RECT 5.330 44.825 1594.550 47.655 ;
        RECT 5.330 39.385 1594.550 42.215 ;
        RECT 5.330 33.945 1594.550 36.775 ;
        RECT 5.330 28.505 1594.550 31.335 ;
        RECT 5.330 23.065 1594.550 25.895 ;
        RECT 5.330 17.625 1594.550 20.455 ;
        RECT 5.330 12.185 1594.550 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1594.360 486.965 ;
      LAYER met1 ;
        RECT 5.520 1.740 1596.590 487.120 ;
      LAYER met2 ;
        RECT 21.070 4.280 1596.560 494.205 ;
        RECT 21.070 1.710 26.490 4.280 ;
        RECT 27.330 1.710 48.570 4.280 ;
        RECT 49.410 1.710 70.650 4.280 ;
        RECT 71.490 1.710 92.730 4.280 ;
        RECT 93.570 1.710 114.810 4.280 ;
        RECT 115.650 1.710 136.890 4.280 ;
        RECT 137.730 1.710 158.970 4.280 ;
        RECT 159.810 1.710 181.050 4.280 ;
        RECT 181.890 1.710 203.130 4.280 ;
        RECT 203.970 1.710 225.210 4.280 ;
        RECT 226.050 1.710 247.290 4.280 ;
        RECT 248.130 1.710 269.370 4.280 ;
        RECT 270.210 1.710 291.450 4.280 ;
        RECT 292.290 1.710 313.530 4.280 ;
        RECT 314.370 1.710 335.610 4.280 ;
        RECT 336.450 1.710 357.690 4.280 ;
        RECT 358.530 1.710 379.770 4.280 ;
        RECT 380.610 1.710 401.850 4.280 ;
        RECT 402.690 1.710 423.930 4.280 ;
        RECT 424.770 1.710 446.010 4.280 ;
        RECT 446.850 1.710 468.090 4.280 ;
        RECT 468.930 1.710 490.170 4.280 ;
        RECT 491.010 1.710 512.250 4.280 ;
        RECT 513.090 1.710 534.330 4.280 ;
        RECT 535.170 1.710 556.410 4.280 ;
        RECT 557.250 1.710 578.490 4.280 ;
        RECT 579.330 1.710 600.570 4.280 ;
        RECT 601.410 1.710 622.650 4.280 ;
        RECT 623.490 1.710 644.730 4.280 ;
        RECT 645.570 1.710 666.810 4.280 ;
        RECT 667.650 1.710 688.890 4.280 ;
        RECT 689.730 1.710 710.970 4.280 ;
        RECT 711.810 1.710 733.050 4.280 ;
        RECT 733.890 1.710 755.130 4.280 ;
        RECT 755.970 1.710 777.210 4.280 ;
        RECT 778.050 1.710 799.290 4.280 ;
        RECT 800.130 1.710 821.370 4.280 ;
        RECT 822.210 1.710 843.450 4.280 ;
        RECT 844.290 1.710 865.530 4.280 ;
        RECT 866.370 1.710 887.610 4.280 ;
        RECT 888.450 1.710 909.690 4.280 ;
        RECT 910.530 1.710 931.770 4.280 ;
        RECT 932.610 1.710 953.850 4.280 ;
        RECT 954.690 1.710 975.930 4.280 ;
        RECT 976.770 1.710 998.010 4.280 ;
        RECT 998.850 1.710 1020.090 4.280 ;
        RECT 1020.930 1.710 1042.170 4.280 ;
        RECT 1043.010 1.710 1064.250 4.280 ;
        RECT 1065.090 1.710 1086.330 4.280 ;
        RECT 1087.170 1.710 1108.410 4.280 ;
        RECT 1109.250 1.710 1130.490 4.280 ;
        RECT 1131.330 1.710 1152.570 4.280 ;
        RECT 1153.410 1.710 1174.650 4.280 ;
        RECT 1175.490 1.710 1196.730 4.280 ;
        RECT 1197.570 1.710 1218.810 4.280 ;
        RECT 1219.650 1.710 1240.890 4.280 ;
        RECT 1241.730 1.710 1262.970 4.280 ;
        RECT 1263.810 1.710 1285.050 4.280 ;
        RECT 1285.890 1.710 1307.130 4.280 ;
        RECT 1307.970 1.710 1329.210 4.280 ;
        RECT 1330.050 1.710 1351.290 4.280 ;
        RECT 1352.130 1.710 1373.370 4.280 ;
        RECT 1374.210 1.710 1395.450 4.280 ;
        RECT 1396.290 1.710 1417.530 4.280 ;
        RECT 1418.370 1.710 1439.610 4.280 ;
        RECT 1440.450 1.710 1461.690 4.280 ;
        RECT 1462.530 1.710 1483.770 4.280 ;
        RECT 1484.610 1.710 1505.850 4.280 ;
        RECT 1506.690 1.710 1527.930 4.280 ;
        RECT 1528.770 1.710 1550.010 4.280 ;
        RECT 1550.850 1.710 1572.090 4.280 ;
        RECT 1572.930 1.710 1596.560 4.280 ;
      LAYER met3 ;
        RECT 21.050 493.320 1595.600 494.185 ;
        RECT 21.050 483.840 1596.135 493.320 ;
        RECT 21.050 482.440 1595.600 483.840 ;
        RECT 21.050 472.960 1596.135 482.440 ;
        RECT 21.050 471.560 1595.600 472.960 ;
        RECT 21.050 462.080 1596.135 471.560 ;
        RECT 21.050 460.680 1595.600 462.080 ;
        RECT 21.050 451.200 1596.135 460.680 ;
        RECT 21.050 449.800 1595.600 451.200 ;
        RECT 21.050 440.320 1596.135 449.800 ;
        RECT 21.050 438.920 1595.600 440.320 ;
        RECT 21.050 429.440 1596.135 438.920 ;
        RECT 21.050 428.040 1595.600 429.440 ;
        RECT 21.050 418.560 1596.135 428.040 ;
        RECT 21.050 417.160 1595.600 418.560 ;
        RECT 21.050 407.680 1596.135 417.160 ;
        RECT 21.050 406.280 1595.600 407.680 ;
        RECT 21.050 396.800 1596.135 406.280 ;
        RECT 21.050 395.400 1595.600 396.800 ;
        RECT 21.050 385.920 1596.135 395.400 ;
        RECT 21.050 384.520 1595.600 385.920 ;
        RECT 21.050 375.040 1596.135 384.520 ;
        RECT 21.050 373.640 1595.600 375.040 ;
        RECT 21.050 364.160 1596.135 373.640 ;
        RECT 21.050 362.760 1595.600 364.160 ;
        RECT 21.050 353.280 1596.135 362.760 ;
        RECT 21.050 351.880 1595.600 353.280 ;
        RECT 21.050 342.400 1596.135 351.880 ;
        RECT 21.050 341.000 1595.600 342.400 ;
        RECT 21.050 331.520 1596.135 341.000 ;
        RECT 21.050 330.120 1595.600 331.520 ;
        RECT 21.050 320.640 1596.135 330.120 ;
        RECT 21.050 319.240 1595.600 320.640 ;
        RECT 21.050 309.760 1596.135 319.240 ;
        RECT 21.050 308.360 1595.600 309.760 ;
        RECT 21.050 298.880 1596.135 308.360 ;
        RECT 21.050 297.480 1595.600 298.880 ;
        RECT 21.050 288.000 1596.135 297.480 ;
        RECT 21.050 286.600 1595.600 288.000 ;
        RECT 21.050 277.120 1596.135 286.600 ;
        RECT 21.050 275.720 1595.600 277.120 ;
        RECT 21.050 266.240 1596.135 275.720 ;
        RECT 21.050 264.840 1595.600 266.240 ;
        RECT 21.050 255.360 1596.135 264.840 ;
        RECT 21.050 253.960 1595.600 255.360 ;
        RECT 21.050 244.480 1596.135 253.960 ;
        RECT 21.050 243.080 1595.600 244.480 ;
        RECT 21.050 233.600 1596.135 243.080 ;
        RECT 21.050 232.200 1595.600 233.600 ;
        RECT 21.050 222.720 1596.135 232.200 ;
        RECT 21.050 221.320 1595.600 222.720 ;
        RECT 21.050 211.840 1596.135 221.320 ;
        RECT 21.050 210.440 1595.600 211.840 ;
        RECT 21.050 200.960 1596.135 210.440 ;
        RECT 21.050 199.560 1595.600 200.960 ;
        RECT 21.050 190.080 1596.135 199.560 ;
        RECT 21.050 188.680 1595.600 190.080 ;
        RECT 21.050 179.200 1596.135 188.680 ;
        RECT 21.050 177.800 1595.600 179.200 ;
        RECT 21.050 168.320 1596.135 177.800 ;
        RECT 21.050 166.920 1595.600 168.320 ;
        RECT 21.050 157.440 1596.135 166.920 ;
        RECT 21.050 156.040 1595.600 157.440 ;
        RECT 21.050 146.560 1596.135 156.040 ;
        RECT 21.050 145.160 1595.600 146.560 ;
        RECT 21.050 135.680 1596.135 145.160 ;
        RECT 21.050 134.280 1595.600 135.680 ;
        RECT 21.050 124.800 1596.135 134.280 ;
        RECT 21.050 123.400 1595.600 124.800 ;
        RECT 21.050 113.920 1596.135 123.400 ;
        RECT 21.050 112.520 1595.600 113.920 ;
        RECT 21.050 103.040 1596.135 112.520 ;
        RECT 21.050 101.640 1595.600 103.040 ;
        RECT 21.050 92.160 1596.135 101.640 ;
        RECT 21.050 90.760 1595.600 92.160 ;
        RECT 21.050 81.280 1596.135 90.760 ;
        RECT 21.050 79.880 1595.600 81.280 ;
        RECT 21.050 70.400 1596.135 79.880 ;
        RECT 21.050 69.000 1595.600 70.400 ;
        RECT 21.050 59.520 1596.135 69.000 ;
        RECT 21.050 58.120 1595.600 59.520 ;
        RECT 21.050 48.640 1596.135 58.120 ;
        RECT 21.050 47.240 1595.600 48.640 ;
        RECT 21.050 37.760 1596.135 47.240 ;
        RECT 21.050 36.360 1595.600 37.760 ;
        RECT 21.050 26.880 1596.135 36.360 ;
        RECT 21.050 25.480 1595.600 26.880 ;
        RECT 21.050 16.000 1596.135 25.480 ;
        RECT 21.050 14.600 1595.600 16.000 ;
        RECT 21.050 5.120 1596.135 14.600 ;
        RECT 21.050 3.720 1595.600 5.120 ;
        RECT 21.050 2.220 1596.135 3.720 ;
      LAYER met4 ;
        RECT 364.615 10.240 404.640 486.025 ;
        RECT 407.040 10.240 481.440 486.025 ;
        RECT 483.840 10.240 558.240 486.025 ;
        RECT 560.640 10.240 635.040 486.025 ;
        RECT 637.440 10.240 711.840 486.025 ;
        RECT 714.240 10.240 788.640 486.025 ;
        RECT 791.040 10.240 865.440 486.025 ;
        RECT 867.840 10.240 942.240 486.025 ;
        RECT 944.640 10.240 1019.040 486.025 ;
        RECT 1021.440 10.240 1095.840 486.025 ;
        RECT 1098.240 10.240 1172.640 486.025 ;
        RECT 1175.040 10.240 1249.440 486.025 ;
        RECT 1251.840 10.240 1326.240 486.025 ;
        RECT 1328.640 10.240 1403.040 486.025 ;
        RECT 1405.440 10.240 1479.840 486.025 ;
        RECT 1482.240 10.240 1556.640 486.025 ;
        RECT 1559.040 10.240 1579.345 486.025 ;
        RECT 364.615 2.215 1579.345 10.240 ;
  END
END SLRV
END LIBRARY

