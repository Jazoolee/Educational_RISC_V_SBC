magic
tech sky130A
magscale 1 2
timestamp 1729343289
<< nwell >>
rect 1066 47045 318910 47366
rect 1066 45957 318910 46523
rect 1066 44869 318910 45435
rect 1066 43781 318910 44347
rect 1066 42693 318910 43259
rect 1066 41605 318910 42171
rect 1066 40517 318910 41083
rect 1066 39429 318910 39995
rect 1066 38341 318910 38907
rect 1066 37253 318910 37819
rect 1066 36165 318910 36731
rect 1066 35077 318910 35643
rect 1066 33989 318910 34555
rect 1066 32901 318910 33467
rect 1066 31813 318910 32379
rect 1066 30725 318910 31291
rect 1066 29637 318910 30203
rect 1066 28549 318910 29115
rect 1066 27461 318910 28027
rect 1066 26373 318910 26939
rect 1066 25285 318910 25851
rect 1066 24197 318910 24763
rect 1066 23109 318910 23675
rect 1066 22021 318910 22587
rect 1066 20933 318910 21499
rect 1066 19845 318910 20411
rect 1066 18757 318910 19323
rect 1066 17669 318910 18235
rect 1066 16581 318910 17147
rect 1066 15493 318910 16059
rect 1066 14405 318910 14971
rect 1066 13317 318910 13883
rect 1066 12229 318910 12795
rect 1066 11141 318910 11707
rect 1066 10053 318910 10619
rect 1066 8965 318910 9531
rect 1066 7877 318910 8443
rect 1066 6789 318910 7355
rect 1066 5701 318910 6267
rect 1066 4613 318910 5179
rect 1066 3525 318910 4091
rect 1066 2437 318910 3003
<< obsli1 >>
rect 1104 2159 318872 47345
<< obsm1 >>
rect 1104 8 318872 47376
<< metal2 >>
rect 5262 0 5318 800
rect 7010 0 7066 800
rect 8758 0 8814 800
rect 10506 0 10562 800
rect 12254 0 12310 800
rect 14002 0 14058 800
rect 15750 0 15806 800
rect 17498 0 17554 800
rect 19246 0 19302 800
rect 20994 0 21050 800
rect 22742 0 22798 800
rect 24490 0 24546 800
rect 26238 0 26294 800
rect 27986 0 28042 800
rect 29734 0 29790 800
rect 31482 0 31538 800
rect 33230 0 33286 800
rect 34978 0 35034 800
rect 36726 0 36782 800
rect 38474 0 38530 800
rect 40222 0 40278 800
rect 41970 0 42026 800
rect 43718 0 43774 800
rect 45466 0 45522 800
rect 47214 0 47270 800
rect 48962 0 49018 800
rect 50710 0 50766 800
rect 52458 0 52514 800
rect 54206 0 54262 800
rect 55954 0 56010 800
rect 57702 0 57758 800
rect 59450 0 59506 800
rect 61198 0 61254 800
rect 62946 0 63002 800
rect 64694 0 64750 800
rect 66442 0 66498 800
rect 68190 0 68246 800
rect 69938 0 69994 800
rect 71686 0 71742 800
rect 73434 0 73490 800
rect 75182 0 75238 800
rect 76930 0 76986 800
rect 78678 0 78734 800
rect 80426 0 80482 800
rect 82174 0 82230 800
rect 83922 0 83978 800
rect 85670 0 85726 800
rect 87418 0 87474 800
rect 89166 0 89222 800
rect 90914 0 90970 800
rect 92662 0 92718 800
rect 94410 0 94466 800
rect 96158 0 96214 800
rect 97906 0 97962 800
rect 99654 0 99710 800
rect 101402 0 101458 800
rect 103150 0 103206 800
rect 104898 0 104954 800
rect 106646 0 106702 800
rect 108394 0 108450 800
rect 110142 0 110198 800
rect 111890 0 111946 800
rect 113638 0 113694 800
rect 115386 0 115442 800
rect 117134 0 117190 800
rect 118882 0 118938 800
rect 120630 0 120686 800
rect 122378 0 122434 800
rect 124126 0 124182 800
rect 125874 0 125930 800
rect 127622 0 127678 800
rect 129370 0 129426 800
rect 131118 0 131174 800
rect 132866 0 132922 800
rect 134614 0 134670 800
rect 136362 0 136418 800
rect 138110 0 138166 800
rect 139858 0 139914 800
rect 141606 0 141662 800
rect 143354 0 143410 800
rect 145102 0 145158 800
rect 146850 0 146906 800
rect 148598 0 148654 800
rect 150346 0 150402 800
rect 152094 0 152150 800
rect 153842 0 153898 800
rect 155590 0 155646 800
rect 157338 0 157394 800
rect 159086 0 159142 800
rect 160834 0 160890 800
rect 162582 0 162638 800
rect 164330 0 164386 800
rect 166078 0 166134 800
rect 167826 0 167882 800
rect 169574 0 169630 800
rect 171322 0 171378 800
rect 173070 0 173126 800
rect 174818 0 174874 800
rect 176566 0 176622 800
rect 178314 0 178370 800
rect 180062 0 180118 800
rect 181810 0 181866 800
rect 183558 0 183614 800
rect 185306 0 185362 800
rect 187054 0 187110 800
rect 188802 0 188858 800
rect 190550 0 190606 800
rect 192298 0 192354 800
rect 194046 0 194102 800
rect 195794 0 195850 800
rect 197542 0 197598 800
rect 199290 0 199346 800
rect 201038 0 201094 800
rect 202786 0 202842 800
rect 204534 0 204590 800
rect 206282 0 206338 800
rect 208030 0 208086 800
rect 209778 0 209834 800
rect 211526 0 211582 800
rect 213274 0 213330 800
rect 215022 0 215078 800
rect 216770 0 216826 800
rect 218518 0 218574 800
rect 220266 0 220322 800
rect 222014 0 222070 800
rect 223762 0 223818 800
rect 225510 0 225566 800
rect 227258 0 227314 800
rect 229006 0 229062 800
rect 230754 0 230810 800
rect 232502 0 232558 800
rect 234250 0 234306 800
rect 235998 0 236054 800
rect 237746 0 237802 800
rect 239494 0 239550 800
rect 241242 0 241298 800
rect 242990 0 243046 800
rect 244738 0 244794 800
rect 246486 0 246542 800
rect 248234 0 248290 800
rect 249982 0 250038 800
rect 251730 0 251786 800
rect 253478 0 253534 800
rect 255226 0 255282 800
rect 256974 0 257030 800
rect 258722 0 258778 800
rect 260470 0 260526 800
rect 262218 0 262274 800
rect 263966 0 264022 800
rect 265714 0 265770 800
rect 267462 0 267518 800
rect 269210 0 269266 800
rect 270958 0 271014 800
rect 272706 0 272762 800
rect 274454 0 274510 800
rect 276202 0 276258 800
rect 277950 0 278006 800
rect 279698 0 279754 800
rect 281446 0 281502 800
rect 283194 0 283250 800
rect 284942 0 284998 800
rect 286690 0 286746 800
rect 288438 0 288494 800
rect 290186 0 290242 800
rect 291934 0 291990 800
rect 293682 0 293738 800
rect 295430 0 295486 800
rect 297178 0 297234 800
rect 298926 0 298982 800
rect 300674 0 300730 800
rect 302422 0 302478 800
rect 304170 0 304226 800
rect 305918 0 305974 800
rect 307666 0 307722 800
rect 309414 0 309470 800
rect 311162 0 311218 800
rect 312910 0 312966 800
rect 314658 0 314714 800
<< obsm2 >>
rect 4214 856 317288 47365
rect 4214 2 5206 856
rect 5374 2 6954 856
rect 7122 2 8702 856
rect 8870 2 10450 856
rect 10618 2 12198 856
rect 12366 2 13946 856
rect 14114 2 15694 856
rect 15862 2 17442 856
rect 17610 2 19190 856
rect 19358 2 20938 856
rect 21106 2 22686 856
rect 22854 2 24434 856
rect 24602 2 26182 856
rect 26350 2 27930 856
rect 28098 2 29678 856
rect 29846 2 31426 856
rect 31594 2 33174 856
rect 33342 2 34922 856
rect 35090 2 36670 856
rect 36838 2 38418 856
rect 38586 2 40166 856
rect 40334 2 41914 856
rect 42082 2 43662 856
rect 43830 2 45410 856
rect 45578 2 47158 856
rect 47326 2 48906 856
rect 49074 2 50654 856
rect 50822 2 52402 856
rect 52570 2 54150 856
rect 54318 2 55898 856
rect 56066 2 57646 856
rect 57814 2 59394 856
rect 59562 2 61142 856
rect 61310 2 62890 856
rect 63058 2 64638 856
rect 64806 2 66386 856
rect 66554 2 68134 856
rect 68302 2 69882 856
rect 70050 2 71630 856
rect 71798 2 73378 856
rect 73546 2 75126 856
rect 75294 2 76874 856
rect 77042 2 78622 856
rect 78790 2 80370 856
rect 80538 2 82118 856
rect 82286 2 83866 856
rect 84034 2 85614 856
rect 85782 2 87362 856
rect 87530 2 89110 856
rect 89278 2 90858 856
rect 91026 2 92606 856
rect 92774 2 94354 856
rect 94522 2 96102 856
rect 96270 2 97850 856
rect 98018 2 99598 856
rect 99766 2 101346 856
rect 101514 2 103094 856
rect 103262 2 104842 856
rect 105010 2 106590 856
rect 106758 2 108338 856
rect 108506 2 110086 856
rect 110254 2 111834 856
rect 112002 2 113582 856
rect 113750 2 115330 856
rect 115498 2 117078 856
rect 117246 2 118826 856
rect 118994 2 120574 856
rect 120742 2 122322 856
rect 122490 2 124070 856
rect 124238 2 125818 856
rect 125986 2 127566 856
rect 127734 2 129314 856
rect 129482 2 131062 856
rect 131230 2 132810 856
rect 132978 2 134558 856
rect 134726 2 136306 856
rect 136474 2 138054 856
rect 138222 2 139802 856
rect 139970 2 141550 856
rect 141718 2 143298 856
rect 143466 2 145046 856
rect 145214 2 146794 856
rect 146962 2 148542 856
rect 148710 2 150290 856
rect 150458 2 152038 856
rect 152206 2 153786 856
rect 153954 2 155534 856
rect 155702 2 157282 856
rect 157450 2 159030 856
rect 159198 2 160778 856
rect 160946 2 162526 856
rect 162694 2 164274 856
rect 164442 2 166022 856
rect 166190 2 167770 856
rect 167938 2 169518 856
rect 169686 2 171266 856
rect 171434 2 173014 856
rect 173182 2 174762 856
rect 174930 2 176510 856
rect 176678 2 178258 856
rect 178426 2 180006 856
rect 180174 2 181754 856
rect 181922 2 183502 856
rect 183670 2 185250 856
rect 185418 2 186998 856
rect 187166 2 188746 856
rect 188914 2 190494 856
rect 190662 2 192242 856
rect 192410 2 193990 856
rect 194158 2 195738 856
rect 195906 2 197486 856
rect 197654 2 199234 856
rect 199402 2 200982 856
rect 201150 2 202730 856
rect 202898 2 204478 856
rect 204646 2 206226 856
rect 206394 2 207974 856
rect 208142 2 209722 856
rect 209890 2 211470 856
rect 211638 2 213218 856
rect 213386 2 214966 856
rect 215134 2 216714 856
rect 216882 2 218462 856
rect 218630 2 220210 856
rect 220378 2 221958 856
rect 222126 2 223706 856
rect 223874 2 225454 856
rect 225622 2 227202 856
rect 227370 2 228950 856
rect 229118 2 230698 856
rect 230866 2 232446 856
rect 232614 2 234194 856
rect 234362 2 235942 856
rect 236110 2 237690 856
rect 237858 2 239438 856
rect 239606 2 241186 856
rect 241354 2 242934 856
rect 243102 2 244682 856
rect 244850 2 246430 856
rect 246598 2 248178 856
rect 248346 2 249926 856
rect 250094 2 251674 856
rect 251842 2 253422 856
rect 253590 2 255170 856
rect 255338 2 256918 856
rect 257086 2 258666 856
rect 258834 2 260414 856
rect 260582 2 262162 856
rect 262330 2 263910 856
rect 264078 2 265658 856
rect 265826 2 267406 856
rect 267574 2 269154 856
rect 269322 2 270902 856
rect 271070 2 272650 856
rect 272818 2 274398 856
rect 274566 2 276146 856
rect 276314 2 277894 856
rect 278062 2 279642 856
rect 279810 2 281390 856
rect 281558 2 283138 856
rect 283306 2 284886 856
rect 285054 2 286634 856
rect 286802 2 288382 856
rect 288550 2 290130 856
rect 290298 2 291878 856
rect 292046 2 293626 856
rect 293794 2 295374 856
rect 295542 2 297122 856
rect 297290 2 298870 856
rect 299038 2 300618 856
rect 300786 2 302366 856
rect 302534 2 304114 856
rect 304282 2 305862 856
rect 306030 2 307610 856
rect 307778 2 309358 856
rect 309526 2 311106 856
rect 311274 2 312854 856
rect 313022 2 314602 856
rect 314770 2 317288 856
<< obsm3 >>
rect 4210 35 316467 47361
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
rect 50288 2128 50608 47376
rect 65648 2128 65968 47376
rect 81008 2128 81328 47376
rect 96368 2128 96688 47376
rect 111728 2128 112048 47376
rect 127088 2128 127408 47376
rect 142448 2128 142768 47376
rect 157808 2128 158128 47376
rect 173168 2128 173488 47376
rect 188528 2128 188848 47376
rect 203888 2128 204208 47376
rect 219248 2128 219568 47376
rect 234608 2128 234928 47376
rect 249968 2128 250288 47376
rect 265328 2128 265648 47376
rect 280688 2128 281008 47376
rect 296048 2128 296368 47376
rect 311408 2128 311728 47376
<< obsm4 >>
rect 61515 2048 65568 39949
rect 66048 2048 80928 39949
rect 81408 2048 96288 39949
rect 96768 2048 111648 39949
rect 112128 2048 127008 39949
rect 127488 2048 142368 39949
rect 142848 2048 157728 39949
rect 158208 2048 173088 39949
rect 173568 2048 188448 39949
rect 188928 2048 203808 39949
rect 204288 2048 219168 39949
rect 219648 2048 234528 39949
rect 235008 2048 249888 39949
rect 250368 2048 265248 39949
rect 265728 2048 280608 39949
rect 281088 2048 295968 39949
rect 296448 2048 300781 39949
rect 61515 35 300781 2048
<< labels >>
rlabel metal2 s 8758 0 8814 800 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 la_data_in[10]
port 2 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 la_data_in[11]
port 3 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[12]
port 4 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[13]
port 5 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[14]
port 6 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[15]
port 7 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[16]
port 8 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[17]
port 9 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 la_data_in[18]
port 10 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[19]
port 11 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_data_in[1]
port 12 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[20]
port 13 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[21]
port 14 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[22]
port 15 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[23]
port 16 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_data_in[24]
port 17 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_data_in[25]
port 18 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_data_in[26]
port 19 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[27]
port 20 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_data_in[28]
port 21 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_data_in[29]
port 22 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 la_data_in[2]
port 23 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[30]
port 24 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_data_in[31]
port 25 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_data_in[32]
port 26 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_data_in[33]
port 27 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[34]
port 28 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_data_in[35]
port 29 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[36]
port 30 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[37]
port 31 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[38]
port 32 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[39]
port 33 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[3]
port 34 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_data_in[40]
port 35 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[41]
port 36 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[42]
port 37 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_data_in[43]
port 38 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[44]
port 39 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[45]
port 40 nsew signal input
rlabel metal2 s 169574 0 169630 800 6 la_data_in[46]
port 41 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_data_in[47]
port 42 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 la_data_in[48]
port 43 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[49]
port 44 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[4]
port 45 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_data_in[50]
port 46 nsew signal input
rlabel metal2 s 187054 0 187110 800 6 la_data_in[51]
port 47 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_data_in[52]
port 48 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_data_in[53]
port 49 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_data_in[54]
port 50 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_data_in[55]
port 51 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_data_in[56]
port 52 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[57]
port 53 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_data_in[58]
port 54 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_data_in[59]
port 55 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[5]
port 56 nsew signal input
rlabel metal2 s 218518 0 218574 800 6 la_data_in[60]
port 57 nsew signal input
rlabel metal2 s 222014 0 222070 800 6 la_data_in[61]
port 58 nsew signal input
rlabel metal2 s 225510 0 225566 800 6 la_data_in[62]
port 59 nsew signal input
rlabel metal2 s 229006 0 229062 800 6 la_data_in[63]
port 60 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_data_in[64]
port 61 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[6]
port 62 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[7]
port 63 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[8]
port 64 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[9]
port 65 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 la_data_out[0]
port 66 nsew signal output
rlabel metal2 s 297178 0 297234 800 6 la_data_out[100]
port 67 nsew signal output
rlabel metal2 s 298926 0 298982 800 6 la_data_out[101]
port 68 nsew signal output
rlabel metal2 s 300674 0 300730 800 6 la_data_out[102]
port 69 nsew signal output
rlabel metal2 s 302422 0 302478 800 6 la_data_out[103]
port 70 nsew signal output
rlabel metal2 s 304170 0 304226 800 6 la_data_out[104]
port 71 nsew signal output
rlabel metal2 s 305918 0 305974 800 6 la_data_out[105]
port 72 nsew signal output
rlabel metal2 s 307666 0 307722 800 6 la_data_out[106]
port 73 nsew signal output
rlabel metal2 s 309414 0 309470 800 6 la_data_out[107]
port 74 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 la_data_out[108]
port 75 nsew signal output
rlabel metal2 s 312910 0 312966 800 6 la_data_out[109]
port 76 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 la_data_out[10]
port 77 nsew signal output
rlabel metal2 s 314658 0 314714 800 6 la_data_out[110]
port 78 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[11]
port 79 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[12]
port 80 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[13]
port 81 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_out[14]
port 82 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[15]
port 83 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_data_out[16]
port 84 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[17]
port 85 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[18]
port 86 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 la_data_out[19]
port 87 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 la_data_out[1]
port 88 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[20]
port 89 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[21]
port 90 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[22]
port 91 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[23]
port 92 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 la_data_out[24]
port 93 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[25]
port 94 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 la_data_out[26]
port 95 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[27]
port 96 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[28]
port 97 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 la_data_out[29]
port 98 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 la_data_out[2]
port 99 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 la_data_out[30]
port 100 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[31]
port 101 nsew signal output
rlabel metal2 s 122378 0 122434 800 6 la_data_out[32]
port 102 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 la_data_out[33]
port 103 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[34]
port 104 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[35]
port 105 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[36]
port 106 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[37]
port 107 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[38]
port 108 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 la_data_out[39]
port 109 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 la_data_out[3]
port 110 nsew signal output
rlabel metal2 s 150346 0 150402 800 6 la_data_out[40]
port 111 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[41]
port 112 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[42]
port 113 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[43]
port 114 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[44]
port 115 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[45]
port 116 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[46]
port 117 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[47]
port 118 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[48]
port 119 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[49]
port 120 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 la_data_out[4]
port 121 nsew signal output
rlabel metal2 s 185306 0 185362 800 6 la_data_out[50]
port 122 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 la_data_out[51]
port 123 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 la_data_out[52]
port 124 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 la_data_out[53]
port 125 nsew signal output
rlabel metal2 s 199290 0 199346 800 6 la_data_out[54]
port 126 nsew signal output
rlabel metal2 s 202786 0 202842 800 6 la_data_out[55]
port 127 nsew signal output
rlabel metal2 s 206282 0 206338 800 6 la_data_out[56]
port 128 nsew signal output
rlabel metal2 s 209778 0 209834 800 6 la_data_out[57]
port 129 nsew signal output
rlabel metal2 s 213274 0 213330 800 6 la_data_out[58]
port 130 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 la_data_out[59]
port 131 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[5]
port 132 nsew signal output
rlabel metal2 s 220266 0 220322 800 6 la_data_out[60]
port 133 nsew signal output
rlabel metal2 s 223762 0 223818 800 6 la_data_out[61]
port 134 nsew signal output
rlabel metal2 s 227258 0 227314 800 6 la_data_out[62]
port 135 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[63]
port 136 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 la_data_out[64]
port 137 nsew signal output
rlabel metal2 s 235998 0 236054 800 6 la_data_out[65]
port 138 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[66]
port 139 nsew signal output
rlabel metal2 s 239494 0 239550 800 6 la_data_out[67]
port 140 nsew signal output
rlabel metal2 s 241242 0 241298 800 6 la_data_out[68]
port 141 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[69]
port 142 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 la_data_out[6]
port 143 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 la_data_out[70]
port 144 nsew signal output
rlabel metal2 s 246486 0 246542 800 6 la_data_out[71]
port 145 nsew signal output
rlabel metal2 s 248234 0 248290 800 6 la_data_out[72]
port 146 nsew signal output
rlabel metal2 s 249982 0 250038 800 6 la_data_out[73]
port 147 nsew signal output
rlabel metal2 s 251730 0 251786 800 6 la_data_out[74]
port 148 nsew signal output
rlabel metal2 s 253478 0 253534 800 6 la_data_out[75]
port 149 nsew signal output
rlabel metal2 s 255226 0 255282 800 6 la_data_out[76]
port 150 nsew signal output
rlabel metal2 s 256974 0 257030 800 6 la_data_out[77]
port 151 nsew signal output
rlabel metal2 s 258722 0 258778 800 6 la_data_out[78]
port 152 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[79]
port 153 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[7]
port 154 nsew signal output
rlabel metal2 s 262218 0 262274 800 6 la_data_out[80]
port 155 nsew signal output
rlabel metal2 s 263966 0 264022 800 6 la_data_out[81]
port 156 nsew signal output
rlabel metal2 s 265714 0 265770 800 6 la_data_out[82]
port 157 nsew signal output
rlabel metal2 s 267462 0 267518 800 6 la_data_out[83]
port 158 nsew signal output
rlabel metal2 s 269210 0 269266 800 6 la_data_out[84]
port 159 nsew signal output
rlabel metal2 s 270958 0 271014 800 6 la_data_out[85]
port 160 nsew signal output
rlabel metal2 s 272706 0 272762 800 6 la_data_out[86]
port 161 nsew signal output
rlabel metal2 s 274454 0 274510 800 6 la_data_out[87]
port 162 nsew signal output
rlabel metal2 s 276202 0 276258 800 6 la_data_out[88]
port 163 nsew signal output
rlabel metal2 s 277950 0 278006 800 6 la_data_out[89]
port 164 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[8]
port 165 nsew signal output
rlabel metal2 s 279698 0 279754 800 6 la_data_out[90]
port 166 nsew signal output
rlabel metal2 s 281446 0 281502 800 6 la_data_out[91]
port 167 nsew signal output
rlabel metal2 s 283194 0 283250 800 6 la_data_out[92]
port 168 nsew signal output
rlabel metal2 s 284942 0 284998 800 6 la_data_out[93]
port 169 nsew signal output
rlabel metal2 s 286690 0 286746 800 6 la_data_out[94]
port 170 nsew signal output
rlabel metal2 s 288438 0 288494 800 6 la_data_out[95]
port 171 nsew signal output
rlabel metal2 s 290186 0 290242 800 6 la_data_out[96]
port 172 nsew signal output
rlabel metal2 s 291934 0 291990 800 6 la_data_out[97]
port 173 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[98]
port 174 nsew signal output
rlabel metal2 s 295430 0 295486 800 6 la_data_out[99]
port 175 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[9]
port 176 nsew signal output
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 47376 6 vccd1
port 177 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 47376 6 vssd1
port 178 nsew ground bidirectional
rlabel metal2 s 5262 0 5318 800 6 wb_clk_i
port 179 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wb_rst_i
port 180 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 320000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 36206410
string GDS_FILE /home/jazoolee/uniccass_example/openlane/user_proj_example/runs/24_10_19_17_54/results/signoff/user_proj_example.magic.gds
string GDS_START 1174994
<< end >>

