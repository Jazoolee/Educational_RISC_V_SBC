magic
tech sky130A
magscale 1 2
timestamp 1730412818
<< nwell >>
rect 1066 80773 256902 81339
rect 1066 79685 256902 80251
rect 1066 78597 256902 79163
rect 1066 77509 256902 78075
rect 1066 76421 256902 76987
rect 1066 75333 256902 75899
rect 1066 74245 256902 74811
rect 1066 73157 256902 73723
rect 1066 72069 256902 72635
rect 1066 70981 256902 71547
rect 1066 69893 256902 70459
rect 1066 68805 256902 69371
rect 1066 67717 256902 68283
rect 1066 66629 256902 67195
rect 1066 65541 256902 66107
rect 1066 64453 256902 65019
rect 1066 63365 256902 63931
rect 1066 62277 256902 62843
rect 1066 61189 256902 61755
rect 1066 60101 256902 60667
rect 1066 59013 256902 59579
rect 1066 57925 256902 58491
rect 1066 56837 256902 57403
rect 1066 55749 256902 56315
rect 1066 54661 256902 55227
rect 1066 53573 256902 54139
rect 1066 52485 256902 53051
rect 1066 51397 256902 51963
rect 1066 50309 256902 50875
rect 1066 49221 256902 49787
rect 1066 48133 256902 48699
rect 1066 47045 256902 47611
rect 1066 45957 256902 46523
rect 1066 44869 256902 45435
rect 1066 43781 256902 44347
rect 1066 42693 256902 43259
rect 1066 41605 256902 42171
rect 1066 40517 256902 41083
rect 1066 39429 256902 39995
rect 1066 38341 256902 38907
rect 1066 37253 256902 37819
rect 1066 36165 256902 36731
rect 1066 35077 256902 35643
rect 1066 33989 256902 34555
rect 1066 32901 256902 33467
rect 1066 31813 256902 32379
rect 1066 30725 256902 31291
rect 1066 29637 256902 30203
rect 1066 28549 256902 29115
rect 1066 27461 256902 28027
rect 1066 26373 256902 26939
rect 1066 25285 256902 25851
rect 1066 24197 256902 24763
rect 1066 23109 256902 23675
rect 1066 22021 256902 22587
rect 1066 20933 256902 21499
rect 1066 19845 256902 20411
rect 1066 18757 256902 19323
rect 1066 17669 256902 18235
rect 1066 16581 256902 17147
rect 1066 15493 256902 16059
rect 1066 14405 256902 14971
rect 1066 13317 256902 13883
rect 1066 12229 256902 12795
rect 1066 11141 256902 11707
rect 1066 10053 256902 10619
rect 1066 8965 256902 9531
rect 1066 7877 256902 8443
rect 1066 6789 256902 7355
rect 1066 5701 256902 6267
rect 1066 4613 256902 5179
rect 1066 3525 256902 4091
rect 1066 2437 256902 3003
<< obsli1 >>
rect 1104 2159 256864 81617
<< obsm1 >>
rect 1104 688 257218 81648
<< metal2 >>
rect 3330 0 3386 800
rect 6918 0 6974 800
rect 10506 0 10562 800
rect 14094 0 14150 800
rect 17682 0 17738 800
rect 21270 0 21326 800
rect 24858 0 24914 800
rect 28446 0 28502 800
rect 32034 0 32090 800
rect 35622 0 35678 800
rect 39210 0 39266 800
rect 42798 0 42854 800
rect 46386 0 46442 800
rect 49974 0 50030 800
rect 53562 0 53618 800
rect 57150 0 57206 800
rect 60738 0 60794 800
rect 64326 0 64382 800
rect 67914 0 67970 800
rect 71502 0 71558 800
rect 75090 0 75146 800
rect 78678 0 78734 800
rect 82266 0 82322 800
rect 85854 0 85910 800
rect 89442 0 89498 800
rect 93030 0 93086 800
rect 96618 0 96674 800
rect 100206 0 100262 800
rect 103794 0 103850 800
rect 107382 0 107438 800
rect 110970 0 111026 800
rect 114558 0 114614 800
rect 118146 0 118202 800
rect 121734 0 121790 800
rect 125322 0 125378 800
rect 128910 0 128966 800
rect 132498 0 132554 800
rect 136086 0 136142 800
rect 139674 0 139730 800
rect 143262 0 143318 800
rect 146850 0 146906 800
rect 150438 0 150494 800
rect 154026 0 154082 800
rect 157614 0 157670 800
rect 161202 0 161258 800
rect 164790 0 164846 800
rect 168378 0 168434 800
rect 171966 0 172022 800
rect 175554 0 175610 800
rect 179142 0 179198 800
rect 182730 0 182786 800
rect 186318 0 186374 800
rect 189906 0 189962 800
rect 193494 0 193550 800
rect 197082 0 197138 800
rect 200670 0 200726 800
rect 204258 0 204314 800
rect 207846 0 207902 800
rect 211434 0 211490 800
rect 215022 0 215078 800
rect 218610 0 218666 800
rect 222198 0 222254 800
rect 225786 0 225842 800
rect 229374 0 229430 800
rect 232962 0 233018 800
rect 236550 0 236606 800
rect 240138 0 240194 800
rect 243726 0 243782 800
rect 247314 0 247370 800
rect 250902 0 250958 800
rect 254490 0 254546 800
<< obsm2 >>
rect 3332 856 257212 81637
rect 3442 575 6862 856
rect 7030 575 10450 856
rect 10618 575 14038 856
rect 14206 575 17626 856
rect 17794 575 21214 856
rect 21382 575 24802 856
rect 24970 575 28390 856
rect 28558 575 31978 856
rect 32146 575 35566 856
rect 35734 575 39154 856
rect 39322 575 42742 856
rect 42910 575 46330 856
rect 46498 575 49918 856
rect 50086 575 53506 856
rect 53674 575 57094 856
rect 57262 575 60682 856
rect 60850 575 64270 856
rect 64438 575 67858 856
rect 68026 575 71446 856
rect 71614 575 75034 856
rect 75202 575 78622 856
rect 78790 575 82210 856
rect 82378 575 85798 856
rect 85966 575 89386 856
rect 89554 575 92974 856
rect 93142 575 96562 856
rect 96730 575 100150 856
rect 100318 575 103738 856
rect 103906 575 107326 856
rect 107494 575 110914 856
rect 111082 575 114502 856
rect 114670 575 118090 856
rect 118258 575 121678 856
rect 121846 575 125266 856
rect 125434 575 128854 856
rect 129022 575 132442 856
rect 132610 575 136030 856
rect 136198 575 139618 856
rect 139786 575 143206 856
rect 143374 575 146794 856
rect 146962 575 150382 856
rect 150550 575 153970 856
rect 154138 575 157558 856
rect 157726 575 161146 856
rect 161314 575 164734 856
rect 164902 575 168322 856
rect 168490 575 171910 856
rect 172078 575 175498 856
rect 175666 575 179086 856
rect 179254 575 182674 856
rect 182842 575 186262 856
rect 186430 575 189850 856
rect 190018 575 193438 856
rect 193606 575 197026 856
rect 197194 575 200614 856
rect 200782 575 204202 856
rect 204370 575 207790 856
rect 207958 575 211378 856
rect 211546 575 214966 856
rect 215134 575 218554 856
rect 218722 575 222142 856
rect 222310 575 225730 856
rect 225898 575 229318 856
rect 229486 575 232906 856
rect 233074 575 236494 856
rect 236662 575 240082 856
rect 240250 575 243670 856
rect 243838 575 247258 856
rect 247426 575 250846 856
rect 251014 575 254434 856
rect 254602 575 257212 856
<< metal3 >>
rect 257200 78616 258000 78736
rect 257200 76984 258000 77104
rect 257200 75352 258000 75472
rect 257200 73720 258000 73840
rect 257200 72088 258000 72208
rect 257200 70456 258000 70576
rect 257200 68824 258000 68944
rect 257200 67192 258000 67312
rect 257200 65560 258000 65680
rect 257200 63928 258000 64048
rect 257200 62296 258000 62416
rect 257200 60664 258000 60784
rect 257200 59032 258000 59152
rect 257200 57400 258000 57520
rect 257200 55768 258000 55888
rect 257200 54136 258000 54256
rect 257200 52504 258000 52624
rect 257200 50872 258000 50992
rect 257200 49240 258000 49360
rect 257200 47608 258000 47728
rect 257200 45976 258000 46096
rect 257200 44344 258000 44464
rect 257200 42712 258000 42832
rect 257200 41080 258000 41200
rect 257200 39448 258000 39568
rect 257200 37816 258000 37936
rect 257200 36184 258000 36304
rect 257200 34552 258000 34672
rect 257200 32920 258000 33040
rect 257200 31288 258000 31408
rect 257200 29656 258000 29776
rect 257200 28024 258000 28144
rect 257200 26392 258000 26512
rect 257200 24760 258000 24880
rect 257200 23128 258000 23248
rect 257200 21496 258000 21616
rect 257200 19864 258000 19984
rect 257200 18232 258000 18352
rect 257200 16600 258000 16720
rect 257200 14968 258000 15088
rect 257200 13336 258000 13456
rect 257200 11704 258000 11824
rect 257200 10072 258000 10192
rect 257200 8440 258000 8560
rect 257200 6808 258000 6928
rect 257200 5176 258000 5296
<< obsm3 >>
rect 4210 78816 257200 81633
rect 4210 78536 257120 78816
rect 4210 77184 257200 78536
rect 4210 76904 257120 77184
rect 4210 75552 257200 76904
rect 4210 75272 257120 75552
rect 4210 73920 257200 75272
rect 4210 73640 257120 73920
rect 4210 72288 257200 73640
rect 4210 72008 257120 72288
rect 4210 70656 257200 72008
rect 4210 70376 257120 70656
rect 4210 69024 257200 70376
rect 4210 68744 257120 69024
rect 4210 67392 257200 68744
rect 4210 67112 257120 67392
rect 4210 65760 257200 67112
rect 4210 65480 257120 65760
rect 4210 64128 257200 65480
rect 4210 63848 257120 64128
rect 4210 62496 257200 63848
rect 4210 62216 257120 62496
rect 4210 60864 257200 62216
rect 4210 60584 257120 60864
rect 4210 59232 257200 60584
rect 4210 58952 257120 59232
rect 4210 57600 257200 58952
rect 4210 57320 257120 57600
rect 4210 55968 257200 57320
rect 4210 55688 257120 55968
rect 4210 54336 257200 55688
rect 4210 54056 257120 54336
rect 4210 52704 257200 54056
rect 4210 52424 257120 52704
rect 4210 51072 257200 52424
rect 4210 50792 257120 51072
rect 4210 49440 257200 50792
rect 4210 49160 257120 49440
rect 4210 47808 257200 49160
rect 4210 47528 257120 47808
rect 4210 46176 257200 47528
rect 4210 45896 257120 46176
rect 4210 44544 257200 45896
rect 4210 44264 257120 44544
rect 4210 42912 257200 44264
rect 4210 42632 257120 42912
rect 4210 41280 257200 42632
rect 4210 41000 257120 41280
rect 4210 39648 257200 41000
rect 4210 39368 257120 39648
rect 4210 38016 257200 39368
rect 4210 37736 257120 38016
rect 4210 36384 257200 37736
rect 4210 36104 257120 36384
rect 4210 34752 257200 36104
rect 4210 34472 257120 34752
rect 4210 33120 257200 34472
rect 4210 32840 257120 33120
rect 4210 31488 257200 32840
rect 4210 31208 257120 31488
rect 4210 29856 257200 31208
rect 4210 29576 257120 29856
rect 4210 28224 257200 29576
rect 4210 27944 257120 28224
rect 4210 26592 257200 27944
rect 4210 26312 257120 26592
rect 4210 24960 257200 26312
rect 4210 24680 257120 24960
rect 4210 23328 257200 24680
rect 4210 23048 257120 23328
rect 4210 21696 257200 23048
rect 4210 21416 257120 21696
rect 4210 20064 257200 21416
rect 4210 19784 257120 20064
rect 4210 18432 257200 19784
rect 4210 18152 257120 18432
rect 4210 16800 257200 18152
rect 4210 16520 257120 16800
rect 4210 15168 257200 16520
rect 4210 14888 257120 15168
rect 4210 13536 257200 14888
rect 4210 13256 257120 13536
rect 4210 11904 257200 13256
rect 4210 11624 257120 11904
rect 4210 10272 257200 11624
rect 4210 9992 257120 10272
rect 4210 8640 257200 9992
rect 4210 8360 257120 8640
rect 4210 7008 257200 8360
rect 4210 6728 257120 7008
rect 4210 5376 257200 6728
rect 4210 5096 257120 5376
rect 4210 579 257200 5096
<< metal4 >>
rect 4208 2128 4528 81648
rect 19568 2128 19888 81648
rect 34928 2128 35248 81648
rect 50288 2128 50608 81648
rect 65648 2128 65968 81648
rect 81008 2128 81328 81648
rect 96368 2128 96688 81648
rect 111728 2128 112048 81648
rect 127088 2128 127408 81648
rect 142448 2128 142768 81648
rect 157808 2128 158128 81648
rect 173168 2128 173488 81648
rect 188528 2128 188848 81648
rect 203888 2128 204208 81648
rect 219248 2128 219568 81648
rect 234608 2128 234928 81648
rect 249968 2128 250288 81648
<< obsm4 >>
rect 26555 2048 34848 78029
rect 35328 2048 50208 78029
rect 50688 2048 65568 78029
rect 66048 2048 80928 78029
rect 81408 2048 96288 78029
rect 96768 2048 111648 78029
rect 112128 2048 127008 78029
rect 127488 2048 142368 78029
rect 142848 2048 157728 78029
rect 158208 2048 173088 78029
rect 173568 2048 188448 78029
rect 188928 2048 203808 78029
rect 204288 2048 219168 78029
rect 219648 2048 234528 78029
rect 235008 2048 249888 78029
rect 250368 2048 255333 78029
rect 26555 579 255333 2048
<< labels >>
rlabel metal2 s 136086 0 136142 800 6 a7[0]
port 1 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 a7[10]
port 2 nsew signal output
rlabel metal2 s 175554 0 175610 800 6 a7[11]
port 3 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 a7[12]
port 4 nsew signal output
rlabel metal2 s 182730 0 182786 800 6 a7[13]
port 5 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 a7[14]
port 6 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 a7[15]
port 7 nsew signal output
rlabel metal2 s 193494 0 193550 800 6 a7[16]
port 8 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 a7[17]
port 9 nsew signal output
rlabel metal2 s 200670 0 200726 800 6 a7[18]
port 10 nsew signal output
rlabel metal2 s 204258 0 204314 800 6 a7[19]
port 11 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 a7[1]
port 12 nsew signal output
rlabel metal2 s 207846 0 207902 800 6 a7[20]
port 13 nsew signal output
rlabel metal2 s 211434 0 211490 800 6 a7[21]
port 14 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 a7[22]
port 15 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 a7[23]
port 16 nsew signal output
rlabel metal2 s 222198 0 222254 800 6 a7[24]
port 17 nsew signal output
rlabel metal2 s 225786 0 225842 800 6 a7[25]
port 18 nsew signal output
rlabel metal2 s 229374 0 229430 800 6 a7[26]
port 19 nsew signal output
rlabel metal2 s 232962 0 233018 800 6 a7[27]
port 20 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 a7[28]
port 21 nsew signal output
rlabel metal2 s 240138 0 240194 800 6 a7[29]
port 22 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 a7[2]
port 23 nsew signal output
rlabel metal2 s 243726 0 243782 800 6 a7[30]
port 24 nsew signal output
rlabel metal2 s 247314 0 247370 800 6 a7[31]
port 25 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 a7[3]
port 26 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 a7[4]
port 27 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 a7[5]
port 28 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 a7[6]
port 29 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 a7[7]
port 30 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 a7[8]
port 31 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 a7[9]
port 32 nsew signal output
rlabel metal3 s 257200 5176 258000 5296 6 csb
port 33 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 gp[0]
port 34 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 gp[10]
port 35 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 gp[11]
port 36 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 gp[12]
port 37 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 gp[13]
port 38 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 gp[14]
port 39 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 gp[15]
port 40 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 gp[16]
port 41 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 gp[17]
port 42 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 gp[18]
port 43 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 gp[19]
port 44 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 gp[1]
port 45 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 gp[20]
port 46 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 gp[21]
port 47 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 gp[22]
port 48 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 gp[23]
port 49 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 gp[24]
port 50 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 gp[25]
port 51 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 gp[26]
port 52 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 gp[27]
port 53 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 gp[28]
port 54 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 gp[29]
port 55 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 gp[2]
port 56 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 gp[30]
port 57 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 gp[31]
port 58 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 gp[3]
port 59 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 gp[4]
port 60 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 gp[5]
port 61 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 gp[6]
port 62 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 gp[7]
port 63 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 gp[8]
port 64 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 gp[9]
port 65 nsew signal output
rlabel metal3 s 257200 65560 258000 65680 6 insMemAddr[0]
port 66 nsew signal output
rlabel metal3 s 257200 67192 258000 67312 6 insMemAddr[1]
port 67 nsew signal output
rlabel metal3 s 257200 68824 258000 68944 6 insMemAddr[2]
port 68 nsew signal output
rlabel metal3 s 257200 70456 258000 70576 6 insMemAddr[3]
port 69 nsew signal output
rlabel metal3 s 257200 72088 258000 72208 6 insMemAddr[4]
port 70 nsew signal output
rlabel metal3 s 257200 73720 258000 73840 6 insMemAddr[5]
port 71 nsew signal output
rlabel metal3 s 257200 75352 258000 75472 6 insMemAddr[6]
port 72 nsew signal output
rlabel metal3 s 257200 76984 258000 77104 6 insMemAddr[7]
port 73 nsew signal output
rlabel metal3 s 257200 78616 258000 78736 6 insMemAddr[8]
port 74 nsew signal output
rlabel metal3 s 257200 13336 258000 13456 6 insMemDataIn[0]
port 75 nsew signal input
rlabel metal3 s 257200 29656 258000 29776 6 insMemDataIn[10]
port 76 nsew signal input
rlabel metal3 s 257200 31288 258000 31408 6 insMemDataIn[11]
port 77 nsew signal input
rlabel metal3 s 257200 32920 258000 33040 6 insMemDataIn[12]
port 78 nsew signal input
rlabel metal3 s 257200 34552 258000 34672 6 insMemDataIn[13]
port 79 nsew signal input
rlabel metal3 s 257200 36184 258000 36304 6 insMemDataIn[14]
port 80 nsew signal input
rlabel metal3 s 257200 37816 258000 37936 6 insMemDataIn[15]
port 81 nsew signal input
rlabel metal3 s 257200 39448 258000 39568 6 insMemDataIn[16]
port 82 nsew signal input
rlabel metal3 s 257200 41080 258000 41200 6 insMemDataIn[17]
port 83 nsew signal input
rlabel metal3 s 257200 42712 258000 42832 6 insMemDataIn[18]
port 84 nsew signal input
rlabel metal3 s 257200 44344 258000 44464 6 insMemDataIn[19]
port 85 nsew signal input
rlabel metal3 s 257200 14968 258000 15088 6 insMemDataIn[1]
port 86 nsew signal input
rlabel metal3 s 257200 45976 258000 46096 6 insMemDataIn[20]
port 87 nsew signal input
rlabel metal3 s 257200 47608 258000 47728 6 insMemDataIn[21]
port 88 nsew signal input
rlabel metal3 s 257200 49240 258000 49360 6 insMemDataIn[22]
port 89 nsew signal input
rlabel metal3 s 257200 50872 258000 50992 6 insMemDataIn[23]
port 90 nsew signal input
rlabel metal3 s 257200 52504 258000 52624 6 insMemDataIn[24]
port 91 nsew signal input
rlabel metal3 s 257200 54136 258000 54256 6 insMemDataIn[25]
port 92 nsew signal input
rlabel metal3 s 257200 55768 258000 55888 6 insMemDataIn[26]
port 93 nsew signal input
rlabel metal3 s 257200 57400 258000 57520 6 insMemDataIn[27]
port 94 nsew signal input
rlabel metal3 s 257200 59032 258000 59152 6 insMemDataIn[28]
port 95 nsew signal input
rlabel metal3 s 257200 60664 258000 60784 6 insMemDataIn[29]
port 96 nsew signal input
rlabel metal3 s 257200 16600 258000 16720 6 insMemDataIn[2]
port 97 nsew signal input
rlabel metal3 s 257200 62296 258000 62416 6 insMemDataIn[30]
port 98 nsew signal input
rlabel metal3 s 257200 63928 258000 64048 6 insMemDataIn[31]
port 99 nsew signal input
rlabel metal3 s 257200 18232 258000 18352 6 insMemDataIn[3]
port 100 nsew signal input
rlabel metal3 s 257200 19864 258000 19984 6 insMemDataIn[4]
port 101 nsew signal input
rlabel metal3 s 257200 21496 258000 21616 6 insMemDataIn[5]
port 102 nsew signal input
rlabel metal3 s 257200 23128 258000 23248 6 insMemDataIn[6]
port 103 nsew signal input
rlabel metal3 s 257200 24760 258000 24880 6 insMemDataIn[7]
port 104 nsew signal input
rlabel metal3 s 257200 26392 258000 26512 6 insMemDataIn[8]
port 105 nsew signal input
rlabel metal3 s 257200 28024 258000 28144 6 insMemDataIn[9]
port 106 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 insMemEn
port 107 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 la_data_in[0]
port 108 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 la_data_in[1]
port 109 nsew signal input
rlabel metal2 s 250902 0 250958 800 6 pc_led
port 110 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 pc_led_oeb
port 111 nsew signal output
rlabel metal4 s 4208 2128 4528 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 81648 6 vccd1
port 112 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 81648 6 vssd1
port 113 nsew ground bidirectional
rlabel metal2 s 3330 0 3386 800 6 wb_clk_i
port 114 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wb_rst_i
port 115 nsew signal input
rlabel metal3 s 257200 6808 258000 6928 6 wmask[0]
port 116 nsew signal output
rlabel metal3 s 257200 8440 258000 8560 6 wmask[1]
port 117 nsew signal output
rlabel metal3 s 257200 10072 258000 10192 6 wmask[2]
port 118 nsew signal output
rlabel metal3 s 257200 11704 258000 11824 6 wmask[3]
port 119 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 258000 84000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 62878988
string GDS_FILE /home/jazoolee/uniccass_example/openlane/SLRV/runs/24_10_31_23_09/results/signoff/SLRV.magic.gds
string GDS_START 1650940
<< end >>

