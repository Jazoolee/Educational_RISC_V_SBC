// This is the unpowered netlist.
module dmem (clock,
    dataMemWen,
    dataMemAddr,
    dataMemDataM2P,
    dataMemDataP2M);
 input clock;
 input dataMemWen;
 input [4:0] dataMemAddr;
 output [31:0] dataMemDataM2P;
 input [31:0] dataMemDataP2M;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire \dataMemory[0][0] ;
 wire \dataMemory[0][10] ;
 wire \dataMemory[0][11] ;
 wire \dataMemory[0][12] ;
 wire \dataMemory[0][13] ;
 wire \dataMemory[0][14] ;
 wire \dataMemory[0][15] ;
 wire \dataMemory[0][16] ;
 wire \dataMemory[0][17] ;
 wire \dataMemory[0][18] ;
 wire \dataMemory[0][19] ;
 wire \dataMemory[0][1] ;
 wire \dataMemory[0][20] ;
 wire \dataMemory[0][21] ;
 wire \dataMemory[0][22] ;
 wire \dataMemory[0][23] ;
 wire \dataMemory[0][24] ;
 wire \dataMemory[0][25] ;
 wire \dataMemory[0][26] ;
 wire \dataMemory[0][27] ;
 wire \dataMemory[0][28] ;
 wire \dataMemory[0][29] ;
 wire \dataMemory[0][2] ;
 wire \dataMemory[0][30] ;
 wire \dataMemory[0][31] ;
 wire \dataMemory[0][3] ;
 wire \dataMemory[0][4] ;
 wire \dataMemory[0][5] ;
 wire \dataMemory[0][6] ;
 wire \dataMemory[0][7] ;
 wire \dataMemory[0][8] ;
 wire \dataMemory[0][9] ;
 wire \dataMemory[10][0] ;
 wire \dataMemory[10][10] ;
 wire \dataMemory[10][11] ;
 wire \dataMemory[10][12] ;
 wire \dataMemory[10][13] ;
 wire \dataMemory[10][14] ;
 wire \dataMemory[10][15] ;
 wire \dataMemory[10][16] ;
 wire \dataMemory[10][17] ;
 wire \dataMemory[10][18] ;
 wire \dataMemory[10][19] ;
 wire \dataMemory[10][1] ;
 wire \dataMemory[10][20] ;
 wire \dataMemory[10][21] ;
 wire \dataMemory[10][22] ;
 wire \dataMemory[10][23] ;
 wire \dataMemory[10][24] ;
 wire \dataMemory[10][25] ;
 wire \dataMemory[10][26] ;
 wire \dataMemory[10][27] ;
 wire \dataMemory[10][28] ;
 wire \dataMemory[10][29] ;
 wire \dataMemory[10][2] ;
 wire \dataMemory[10][30] ;
 wire \dataMemory[10][31] ;
 wire \dataMemory[10][3] ;
 wire \dataMemory[10][4] ;
 wire \dataMemory[10][5] ;
 wire \dataMemory[10][6] ;
 wire \dataMemory[10][7] ;
 wire \dataMemory[10][8] ;
 wire \dataMemory[10][9] ;
 wire \dataMemory[11][0] ;
 wire \dataMemory[11][10] ;
 wire \dataMemory[11][11] ;
 wire \dataMemory[11][12] ;
 wire \dataMemory[11][13] ;
 wire \dataMemory[11][14] ;
 wire \dataMemory[11][15] ;
 wire \dataMemory[11][16] ;
 wire \dataMemory[11][17] ;
 wire \dataMemory[11][18] ;
 wire \dataMemory[11][19] ;
 wire \dataMemory[11][1] ;
 wire \dataMemory[11][20] ;
 wire \dataMemory[11][21] ;
 wire \dataMemory[11][22] ;
 wire \dataMemory[11][23] ;
 wire \dataMemory[11][24] ;
 wire \dataMemory[11][25] ;
 wire \dataMemory[11][26] ;
 wire \dataMemory[11][27] ;
 wire \dataMemory[11][28] ;
 wire \dataMemory[11][29] ;
 wire \dataMemory[11][2] ;
 wire \dataMemory[11][30] ;
 wire \dataMemory[11][31] ;
 wire \dataMemory[11][3] ;
 wire \dataMemory[11][4] ;
 wire \dataMemory[11][5] ;
 wire \dataMemory[11][6] ;
 wire \dataMemory[11][7] ;
 wire \dataMemory[11][8] ;
 wire \dataMemory[11][9] ;
 wire \dataMemory[12][0] ;
 wire \dataMemory[12][10] ;
 wire \dataMemory[12][11] ;
 wire \dataMemory[12][12] ;
 wire \dataMemory[12][13] ;
 wire \dataMemory[12][14] ;
 wire \dataMemory[12][15] ;
 wire \dataMemory[12][16] ;
 wire \dataMemory[12][17] ;
 wire \dataMemory[12][18] ;
 wire \dataMemory[12][19] ;
 wire \dataMemory[12][1] ;
 wire \dataMemory[12][20] ;
 wire \dataMemory[12][21] ;
 wire \dataMemory[12][22] ;
 wire \dataMemory[12][23] ;
 wire \dataMemory[12][24] ;
 wire \dataMemory[12][25] ;
 wire \dataMemory[12][26] ;
 wire \dataMemory[12][27] ;
 wire \dataMemory[12][28] ;
 wire \dataMemory[12][29] ;
 wire \dataMemory[12][2] ;
 wire \dataMemory[12][30] ;
 wire \dataMemory[12][31] ;
 wire \dataMemory[12][3] ;
 wire \dataMemory[12][4] ;
 wire \dataMemory[12][5] ;
 wire \dataMemory[12][6] ;
 wire \dataMemory[12][7] ;
 wire \dataMemory[12][8] ;
 wire \dataMemory[12][9] ;
 wire \dataMemory[13][0] ;
 wire \dataMemory[13][10] ;
 wire \dataMemory[13][11] ;
 wire \dataMemory[13][12] ;
 wire \dataMemory[13][13] ;
 wire \dataMemory[13][14] ;
 wire \dataMemory[13][15] ;
 wire \dataMemory[13][16] ;
 wire \dataMemory[13][17] ;
 wire \dataMemory[13][18] ;
 wire \dataMemory[13][19] ;
 wire \dataMemory[13][1] ;
 wire \dataMemory[13][20] ;
 wire \dataMemory[13][21] ;
 wire \dataMemory[13][22] ;
 wire \dataMemory[13][23] ;
 wire \dataMemory[13][24] ;
 wire \dataMemory[13][25] ;
 wire \dataMemory[13][26] ;
 wire \dataMemory[13][27] ;
 wire \dataMemory[13][28] ;
 wire \dataMemory[13][29] ;
 wire \dataMemory[13][2] ;
 wire \dataMemory[13][30] ;
 wire \dataMemory[13][31] ;
 wire \dataMemory[13][3] ;
 wire \dataMemory[13][4] ;
 wire \dataMemory[13][5] ;
 wire \dataMemory[13][6] ;
 wire \dataMemory[13][7] ;
 wire \dataMemory[13][8] ;
 wire \dataMemory[13][9] ;
 wire \dataMemory[14][0] ;
 wire \dataMemory[14][10] ;
 wire \dataMemory[14][11] ;
 wire \dataMemory[14][12] ;
 wire \dataMemory[14][13] ;
 wire \dataMemory[14][14] ;
 wire \dataMemory[14][15] ;
 wire \dataMemory[14][16] ;
 wire \dataMemory[14][17] ;
 wire \dataMemory[14][18] ;
 wire \dataMemory[14][19] ;
 wire \dataMemory[14][1] ;
 wire \dataMemory[14][20] ;
 wire \dataMemory[14][21] ;
 wire \dataMemory[14][22] ;
 wire \dataMemory[14][23] ;
 wire \dataMemory[14][24] ;
 wire \dataMemory[14][25] ;
 wire \dataMemory[14][26] ;
 wire \dataMemory[14][27] ;
 wire \dataMemory[14][28] ;
 wire \dataMemory[14][29] ;
 wire \dataMemory[14][2] ;
 wire \dataMemory[14][30] ;
 wire \dataMemory[14][31] ;
 wire \dataMemory[14][3] ;
 wire \dataMemory[14][4] ;
 wire \dataMemory[14][5] ;
 wire \dataMemory[14][6] ;
 wire \dataMemory[14][7] ;
 wire \dataMemory[14][8] ;
 wire \dataMemory[14][9] ;
 wire \dataMemory[15][0] ;
 wire \dataMemory[15][10] ;
 wire \dataMemory[15][11] ;
 wire \dataMemory[15][12] ;
 wire \dataMemory[15][13] ;
 wire \dataMemory[15][14] ;
 wire \dataMemory[15][15] ;
 wire \dataMemory[15][16] ;
 wire \dataMemory[15][17] ;
 wire \dataMemory[15][18] ;
 wire \dataMemory[15][19] ;
 wire \dataMemory[15][1] ;
 wire \dataMemory[15][20] ;
 wire \dataMemory[15][21] ;
 wire \dataMemory[15][22] ;
 wire \dataMemory[15][23] ;
 wire \dataMemory[15][24] ;
 wire \dataMemory[15][25] ;
 wire \dataMemory[15][26] ;
 wire \dataMemory[15][27] ;
 wire \dataMemory[15][28] ;
 wire \dataMemory[15][29] ;
 wire \dataMemory[15][2] ;
 wire \dataMemory[15][30] ;
 wire \dataMemory[15][31] ;
 wire \dataMemory[15][3] ;
 wire \dataMemory[15][4] ;
 wire \dataMemory[15][5] ;
 wire \dataMemory[15][6] ;
 wire \dataMemory[15][7] ;
 wire \dataMemory[15][8] ;
 wire \dataMemory[15][9] ;
 wire \dataMemory[16][0] ;
 wire \dataMemory[16][10] ;
 wire \dataMemory[16][11] ;
 wire \dataMemory[16][12] ;
 wire \dataMemory[16][13] ;
 wire \dataMemory[16][14] ;
 wire \dataMemory[16][15] ;
 wire \dataMemory[16][16] ;
 wire \dataMemory[16][17] ;
 wire \dataMemory[16][18] ;
 wire \dataMemory[16][19] ;
 wire \dataMemory[16][1] ;
 wire \dataMemory[16][20] ;
 wire \dataMemory[16][21] ;
 wire \dataMemory[16][22] ;
 wire \dataMemory[16][23] ;
 wire \dataMemory[16][24] ;
 wire \dataMemory[16][25] ;
 wire \dataMemory[16][26] ;
 wire \dataMemory[16][27] ;
 wire \dataMemory[16][28] ;
 wire \dataMemory[16][29] ;
 wire \dataMemory[16][2] ;
 wire \dataMemory[16][30] ;
 wire \dataMemory[16][31] ;
 wire \dataMemory[16][3] ;
 wire \dataMemory[16][4] ;
 wire \dataMemory[16][5] ;
 wire \dataMemory[16][6] ;
 wire \dataMemory[16][7] ;
 wire \dataMemory[16][8] ;
 wire \dataMemory[16][9] ;
 wire \dataMemory[17][0] ;
 wire \dataMemory[17][10] ;
 wire \dataMemory[17][11] ;
 wire \dataMemory[17][12] ;
 wire \dataMemory[17][13] ;
 wire \dataMemory[17][14] ;
 wire \dataMemory[17][15] ;
 wire \dataMemory[17][16] ;
 wire \dataMemory[17][17] ;
 wire \dataMemory[17][18] ;
 wire \dataMemory[17][19] ;
 wire \dataMemory[17][1] ;
 wire \dataMemory[17][20] ;
 wire \dataMemory[17][21] ;
 wire \dataMemory[17][22] ;
 wire \dataMemory[17][23] ;
 wire \dataMemory[17][24] ;
 wire \dataMemory[17][25] ;
 wire \dataMemory[17][26] ;
 wire \dataMemory[17][27] ;
 wire \dataMemory[17][28] ;
 wire \dataMemory[17][29] ;
 wire \dataMemory[17][2] ;
 wire \dataMemory[17][30] ;
 wire \dataMemory[17][31] ;
 wire \dataMemory[17][3] ;
 wire \dataMemory[17][4] ;
 wire \dataMemory[17][5] ;
 wire \dataMemory[17][6] ;
 wire \dataMemory[17][7] ;
 wire \dataMemory[17][8] ;
 wire \dataMemory[17][9] ;
 wire \dataMemory[18][0] ;
 wire \dataMemory[18][10] ;
 wire \dataMemory[18][11] ;
 wire \dataMemory[18][12] ;
 wire \dataMemory[18][13] ;
 wire \dataMemory[18][14] ;
 wire \dataMemory[18][15] ;
 wire \dataMemory[18][16] ;
 wire \dataMemory[18][17] ;
 wire \dataMemory[18][18] ;
 wire \dataMemory[18][19] ;
 wire \dataMemory[18][1] ;
 wire \dataMemory[18][20] ;
 wire \dataMemory[18][21] ;
 wire \dataMemory[18][22] ;
 wire \dataMemory[18][23] ;
 wire \dataMemory[18][24] ;
 wire \dataMemory[18][25] ;
 wire \dataMemory[18][26] ;
 wire \dataMemory[18][27] ;
 wire \dataMemory[18][28] ;
 wire \dataMemory[18][29] ;
 wire \dataMemory[18][2] ;
 wire \dataMemory[18][30] ;
 wire \dataMemory[18][31] ;
 wire \dataMemory[18][3] ;
 wire \dataMemory[18][4] ;
 wire \dataMemory[18][5] ;
 wire \dataMemory[18][6] ;
 wire \dataMemory[18][7] ;
 wire \dataMemory[18][8] ;
 wire \dataMemory[18][9] ;
 wire \dataMemory[19][0] ;
 wire \dataMemory[19][10] ;
 wire \dataMemory[19][11] ;
 wire \dataMemory[19][12] ;
 wire \dataMemory[19][13] ;
 wire \dataMemory[19][14] ;
 wire \dataMemory[19][15] ;
 wire \dataMemory[19][16] ;
 wire \dataMemory[19][17] ;
 wire \dataMemory[19][18] ;
 wire \dataMemory[19][19] ;
 wire \dataMemory[19][1] ;
 wire \dataMemory[19][20] ;
 wire \dataMemory[19][21] ;
 wire \dataMemory[19][22] ;
 wire \dataMemory[19][23] ;
 wire \dataMemory[19][24] ;
 wire \dataMemory[19][25] ;
 wire \dataMemory[19][26] ;
 wire \dataMemory[19][27] ;
 wire \dataMemory[19][28] ;
 wire \dataMemory[19][29] ;
 wire \dataMemory[19][2] ;
 wire \dataMemory[19][30] ;
 wire \dataMemory[19][31] ;
 wire \dataMemory[19][3] ;
 wire \dataMemory[19][4] ;
 wire \dataMemory[19][5] ;
 wire \dataMemory[19][6] ;
 wire \dataMemory[19][7] ;
 wire \dataMemory[19][8] ;
 wire \dataMemory[19][9] ;
 wire \dataMemory[1][0] ;
 wire \dataMemory[1][10] ;
 wire \dataMemory[1][11] ;
 wire \dataMemory[1][12] ;
 wire \dataMemory[1][13] ;
 wire \dataMemory[1][14] ;
 wire \dataMemory[1][15] ;
 wire \dataMemory[1][16] ;
 wire \dataMemory[1][17] ;
 wire \dataMemory[1][18] ;
 wire \dataMemory[1][19] ;
 wire \dataMemory[1][1] ;
 wire \dataMemory[1][20] ;
 wire \dataMemory[1][21] ;
 wire \dataMemory[1][22] ;
 wire \dataMemory[1][23] ;
 wire \dataMemory[1][24] ;
 wire \dataMemory[1][25] ;
 wire \dataMemory[1][26] ;
 wire \dataMemory[1][27] ;
 wire \dataMemory[1][28] ;
 wire \dataMemory[1][29] ;
 wire \dataMemory[1][2] ;
 wire \dataMemory[1][30] ;
 wire \dataMemory[1][31] ;
 wire \dataMemory[1][3] ;
 wire \dataMemory[1][4] ;
 wire \dataMemory[1][5] ;
 wire \dataMemory[1][6] ;
 wire \dataMemory[1][7] ;
 wire \dataMemory[1][8] ;
 wire \dataMemory[1][9] ;
 wire \dataMemory[20][0] ;
 wire \dataMemory[20][10] ;
 wire \dataMemory[20][11] ;
 wire \dataMemory[20][12] ;
 wire \dataMemory[20][13] ;
 wire \dataMemory[20][14] ;
 wire \dataMemory[20][15] ;
 wire \dataMemory[20][16] ;
 wire \dataMemory[20][17] ;
 wire \dataMemory[20][18] ;
 wire \dataMemory[20][19] ;
 wire \dataMemory[20][1] ;
 wire \dataMemory[20][20] ;
 wire \dataMemory[20][21] ;
 wire \dataMemory[20][22] ;
 wire \dataMemory[20][23] ;
 wire \dataMemory[20][24] ;
 wire \dataMemory[20][25] ;
 wire \dataMemory[20][26] ;
 wire \dataMemory[20][27] ;
 wire \dataMemory[20][28] ;
 wire \dataMemory[20][29] ;
 wire \dataMemory[20][2] ;
 wire \dataMemory[20][30] ;
 wire \dataMemory[20][31] ;
 wire \dataMemory[20][3] ;
 wire \dataMemory[20][4] ;
 wire \dataMemory[20][5] ;
 wire \dataMemory[20][6] ;
 wire \dataMemory[20][7] ;
 wire \dataMemory[20][8] ;
 wire \dataMemory[20][9] ;
 wire \dataMemory[21][0] ;
 wire \dataMemory[21][10] ;
 wire \dataMemory[21][11] ;
 wire \dataMemory[21][12] ;
 wire \dataMemory[21][13] ;
 wire \dataMemory[21][14] ;
 wire \dataMemory[21][15] ;
 wire \dataMemory[21][16] ;
 wire \dataMemory[21][17] ;
 wire \dataMemory[21][18] ;
 wire \dataMemory[21][19] ;
 wire \dataMemory[21][1] ;
 wire \dataMemory[21][20] ;
 wire \dataMemory[21][21] ;
 wire \dataMemory[21][22] ;
 wire \dataMemory[21][23] ;
 wire \dataMemory[21][24] ;
 wire \dataMemory[21][25] ;
 wire \dataMemory[21][26] ;
 wire \dataMemory[21][27] ;
 wire \dataMemory[21][28] ;
 wire \dataMemory[21][29] ;
 wire \dataMemory[21][2] ;
 wire \dataMemory[21][30] ;
 wire \dataMemory[21][31] ;
 wire \dataMemory[21][3] ;
 wire \dataMemory[21][4] ;
 wire \dataMemory[21][5] ;
 wire \dataMemory[21][6] ;
 wire \dataMemory[21][7] ;
 wire \dataMemory[21][8] ;
 wire \dataMemory[21][9] ;
 wire \dataMemory[22][0] ;
 wire \dataMemory[22][10] ;
 wire \dataMemory[22][11] ;
 wire \dataMemory[22][12] ;
 wire \dataMemory[22][13] ;
 wire \dataMemory[22][14] ;
 wire \dataMemory[22][15] ;
 wire \dataMemory[22][16] ;
 wire \dataMemory[22][17] ;
 wire \dataMemory[22][18] ;
 wire \dataMemory[22][19] ;
 wire \dataMemory[22][1] ;
 wire \dataMemory[22][20] ;
 wire \dataMemory[22][21] ;
 wire \dataMemory[22][22] ;
 wire \dataMemory[22][23] ;
 wire \dataMemory[22][24] ;
 wire \dataMemory[22][25] ;
 wire \dataMemory[22][26] ;
 wire \dataMemory[22][27] ;
 wire \dataMemory[22][28] ;
 wire \dataMemory[22][29] ;
 wire \dataMemory[22][2] ;
 wire \dataMemory[22][30] ;
 wire \dataMemory[22][31] ;
 wire \dataMemory[22][3] ;
 wire \dataMemory[22][4] ;
 wire \dataMemory[22][5] ;
 wire \dataMemory[22][6] ;
 wire \dataMemory[22][7] ;
 wire \dataMemory[22][8] ;
 wire \dataMemory[22][9] ;
 wire \dataMemory[23][0] ;
 wire \dataMemory[23][10] ;
 wire \dataMemory[23][11] ;
 wire \dataMemory[23][12] ;
 wire \dataMemory[23][13] ;
 wire \dataMemory[23][14] ;
 wire \dataMemory[23][15] ;
 wire \dataMemory[23][16] ;
 wire \dataMemory[23][17] ;
 wire \dataMemory[23][18] ;
 wire \dataMemory[23][19] ;
 wire \dataMemory[23][1] ;
 wire \dataMemory[23][20] ;
 wire \dataMemory[23][21] ;
 wire \dataMemory[23][22] ;
 wire \dataMemory[23][23] ;
 wire \dataMemory[23][24] ;
 wire \dataMemory[23][25] ;
 wire \dataMemory[23][26] ;
 wire \dataMemory[23][27] ;
 wire \dataMemory[23][28] ;
 wire \dataMemory[23][29] ;
 wire \dataMemory[23][2] ;
 wire \dataMemory[23][30] ;
 wire \dataMemory[23][31] ;
 wire \dataMemory[23][3] ;
 wire \dataMemory[23][4] ;
 wire \dataMemory[23][5] ;
 wire \dataMemory[23][6] ;
 wire \dataMemory[23][7] ;
 wire \dataMemory[23][8] ;
 wire \dataMemory[23][9] ;
 wire \dataMemory[24][0] ;
 wire \dataMemory[24][10] ;
 wire \dataMemory[24][11] ;
 wire \dataMemory[24][12] ;
 wire \dataMemory[24][13] ;
 wire \dataMemory[24][14] ;
 wire \dataMemory[24][15] ;
 wire \dataMemory[24][16] ;
 wire \dataMemory[24][17] ;
 wire \dataMemory[24][18] ;
 wire \dataMemory[24][19] ;
 wire \dataMemory[24][1] ;
 wire \dataMemory[24][20] ;
 wire \dataMemory[24][21] ;
 wire \dataMemory[24][22] ;
 wire \dataMemory[24][23] ;
 wire \dataMemory[24][24] ;
 wire \dataMemory[24][25] ;
 wire \dataMemory[24][26] ;
 wire \dataMemory[24][27] ;
 wire \dataMemory[24][28] ;
 wire \dataMemory[24][29] ;
 wire \dataMemory[24][2] ;
 wire \dataMemory[24][30] ;
 wire \dataMemory[24][31] ;
 wire \dataMemory[24][3] ;
 wire \dataMemory[24][4] ;
 wire \dataMemory[24][5] ;
 wire \dataMemory[24][6] ;
 wire \dataMemory[24][7] ;
 wire \dataMemory[24][8] ;
 wire \dataMemory[24][9] ;
 wire \dataMemory[25][0] ;
 wire \dataMemory[25][10] ;
 wire \dataMemory[25][11] ;
 wire \dataMemory[25][12] ;
 wire \dataMemory[25][13] ;
 wire \dataMemory[25][14] ;
 wire \dataMemory[25][15] ;
 wire \dataMemory[25][16] ;
 wire \dataMemory[25][17] ;
 wire \dataMemory[25][18] ;
 wire \dataMemory[25][19] ;
 wire \dataMemory[25][1] ;
 wire \dataMemory[25][20] ;
 wire \dataMemory[25][21] ;
 wire \dataMemory[25][22] ;
 wire \dataMemory[25][23] ;
 wire \dataMemory[25][24] ;
 wire \dataMemory[25][25] ;
 wire \dataMemory[25][26] ;
 wire \dataMemory[25][27] ;
 wire \dataMemory[25][28] ;
 wire \dataMemory[25][29] ;
 wire \dataMemory[25][2] ;
 wire \dataMemory[25][30] ;
 wire \dataMemory[25][31] ;
 wire \dataMemory[25][3] ;
 wire \dataMemory[25][4] ;
 wire \dataMemory[25][5] ;
 wire \dataMemory[25][6] ;
 wire \dataMemory[25][7] ;
 wire \dataMemory[25][8] ;
 wire \dataMemory[25][9] ;
 wire \dataMemory[26][0] ;
 wire \dataMemory[26][10] ;
 wire \dataMemory[26][11] ;
 wire \dataMemory[26][12] ;
 wire \dataMemory[26][13] ;
 wire \dataMemory[26][14] ;
 wire \dataMemory[26][15] ;
 wire \dataMemory[26][16] ;
 wire \dataMemory[26][17] ;
 wire \dataMemory[26][18] ;
 wire \dataMemory[26][19] ;
 wire \dataMemory[26][1] ;
 wire \dataMemory[26][20] ;
 wire \dataMemory[26][21] ;
 wire \dataMemory[26][22] ;
 wire \dataMemory[26][23] ;
 wire \dataMemory[26][24] ;
 wire \dataMemory[26][25] ;
 wire \dataMemory[26][26] ;
 wire \dataMemory[26][27] ;
 wire \dataMemory[26][28] ;
 wire \dataMemory[26][29] ;
 wire \dataMemory[26][2] ;
 wire \dataMemory[26][30] ;
 wire \dataMemory[26][31] ;
 wire \dataMemory[26][3] ;
 wire \dataMemory[26][4] ;
 wire \dataMemory[26][5] ;
 wire \dataMemory[26][6] ;
 wire \dataMemory[26][7] ;
 wire \dataMemory[26][8] ;
 wire \dataMemory[26][9] ;
 wire \dataMemory[27][0] ;
 wire \dataMemory[27][10] ;
 wire \dataMemory[27][11] ;
 wire \dataMemory[27][12] ;
 wire \dataMemory[27][13] ;
 wire \dataMemory[27][14] ;
 wire \dataMemory[27][15] ;
 wire \dataMemory[27][16] ;
 wire \dataMemory[27][17] ;
 wire \dataMemory[27][18] ;
 wire \dataMemory[27][19] ;
 wire \dataMemory[27][1] ;
 wire \dataMemory[27][20] ;
 wire \dataMemory[27][21] ;
 wire \dataMemory[27][22] ;
 wire \dataMemory[27][23] ;
 wire \dataMemory[27][24] ;
 wire \dataMemory[27][25] ;
 wire \dataMemory[27][26] ;
 wire \dataMemory[27][27] ;
 wire \dataMemory[27][28] ;
 wire \dataMemory[27][29] ;
 wire \dataMemory[27][2] ;
 wire \dataMemory[27][30] ;
 wire \dataMemory[27][31] ;
 wire \dataMemory[27][3] ;
 wire \dataMemory[27][4] ;
 wire \dataMemory[27][5] ;
 wire \dataMemory[27][6] ;
 wire \dataMemory[27][7] ;
 wire \dataMemory[27][8] ;
 wire \dataMemory[27][9] ;
 wire \dataMemory[28][0] ;
 wire \dataMemory[28][10] ;
 wire \dataMemory[28][11] ;
 wire \dataMemory[28][12] ;
 wire \dataMemory[28][13] ;
 wire \dataMemory[28][14] ;
 wire \dataMemory[28][15] ;
 wire \dataMemory[28][16] ;
 wire \dataMemory[28][17] ;
 wire \dataMemory[28][18] ;
 wire \dataMemory[28][19] ;
 wire \dataMemory[28][1] ;
 wire \dataMemory[28][20] ;
 wire \dataMemory[28][21] ;
 wire \dataMemory[28][22] ;
 wire \dataMemory[28][23] ;
 wire \dataMemory[28][24] ;
 wire \dataMemory[28][25] ;
 wire \dataMemory[28][26] ;
 wire \dataMemory[28][27] ;
 wire \dataMemory[28][28] ;
 wire \dataMemory[28][29] ;
 wire \dataMemory[28][2] ;
 wire \dataMemory[28][30] ;
 wire \dataMemory[28][31] ;
 wire \dataMemory[28][3] ;
 wire \dataMemory[28][4] ;
 wire \dataMemory[28][5] ;
 wire \dataMemory[28][6] ;
 wire \dataMemory[28][7] ;
 wire \dataMemory[28][8] ;
 wire \dataMemory[28][9] ;
 wire \dataMemory[29][0] ;
 wire \dataMemory[29][10] ;
 wire \dataMemory[29][11] ;
 wire \dataMemory[29][12] ;
 wire \dataMemory[29][13] ;
 wire \dataMemory[29][14] ;
 wire \dataMemory[29][15] ;
 wire \dataMemory[29][16] ;
 wire \dataMemory[29][17] ;
 wire \dataMemory[29][18] ;
 wire \dataMemory[29][19] ;
 wire \dataMemory[29][1] ;
 wire \dataMemory[29][20] ;
 wire \dataMemory[29][21] ;
 wire \dataMemory[29][22] ;
 wire \dataMemory[29][23] ;
 wire \dataMemory[29][24] ;
 wire \dataMemory[29][25] ;
 wire \dataMemory[29][26] ;
 wire \dataMemory[29][27] ;
 wire \dataMemory[29][28] ;
 wire \dataMemory[29][29] ;
 wire \dataMemory[29][2] ;
 wire \dataMemory[29][30] ;
 wire \dataMemory[29][31] ;
 wire \dataMemory[29][3] ;
 wire \dataMemory[29][4] ;
 wire \dataMemory[29][5] ;
 wire \dataMemory[29][6] ;
 wire \dataMemory[29][7] ;
 wire \dataMemory[29][8] ;
 wire \dataMemory[29][9] ;
 wire \dataMemory[2][0] ;
 wire \dataMemory[2][10] ;
 wire \dataMemory[2][11] ;
 wire \dataMemory[2][12] ;
 wire \dataMemory[2][13] ;
 wire \dataMemory[2][14] ;
 wire \dataMemory[2][15] ;
 wire \dataMemory[2][16] ;
 wire \dataMemory[2][17] ;
 wire \dataMemory[2][18] ;
 wire \dataMemory[2][19] ;
 wire \dataMemory[2][1] ;
 wire \dataMemory[2][20] ;
 wire \dataMemory[2][21] ;
 wire \dataMemory[2][22] ;
 wire \dataMemory[2][23] ;
 wire \dataMemory[2][24] ;
 wire \dataMemory[2][25] ;
 wire \dataMemory[2][26] ;
 wire \dataMemory[2][27] ;
 wire \dataMemory[2][28] ;
 wire \dataMemory[2][29] ;
 wire \dataMemory[2][2] ;
 wire \dataMemory[2][30] ;
 wire \dataMemory[2][31] ;
 wire \dataMemory[2][3] ;
 wire \dataMemory[2][4] ;
 wire \dataMemory[2][5] ;
 wire \dataMemory[2][6] ;
 wire \dataMemory[2][7] ;
 wire \dataMemory[2][8] ;
 wire \dataMemory[2][9] ;
 wire \dataMemory[30][0] ;
 wire \dataMemory[30][10] ;
 wire \dataMemory[30][11] ;
 wire \dataMemory[30][12] ;
 wire \dataMemory[30][13] ;
 wire \dataMemory[30][14] ;
 wire \dataMemory[30][15] ;
 wire \dataMemory[30][16] ;
 wire \dataMemory[30][17] ;
 wire \dataMemory[30][18] ;
 wire \dataMemory[30][19] ;
 wire \dataMemory[30][1] ;
 wire \dataMemory[30][20] ;
 wire \dataMemory[30][21] ;
 wire \dataMemory[30][22] ;
 wire \dataMemory[30][23] ;
 wire \dataMemory[30][24] ;
 wire \dataMemory[30][25] ;
 wire \dataMemory[30][26] ;
 wire \dataMemory[30][27] ;
 wire \dataMemory[30][28] ;
 wire \dataMemory[30][29] ;
 wire \dataMemory[30][2] ;
 wire \dataMemory[30][30] ;
 wire \dataMemory[30][31] ;
 wire \dataMemory[30][3] ;
 wire \dataMemory[30][4] ;
 wire \dataMemory[30][5] ;
 wire \dataMemory[30][6] ;
 wire \dataMemory[30][7] ;
 wire \dataMemory[30][8] ;
 wire \dataMemory[30][9] ;
 wire \dataMemory[31][0] ;
 wire \dataMemory[31][10] ;
 wire \dataMemory[31][11] ;
 wire \dataMemory[31][12] ;
 wire \dataMemory[31][13] ;
 wire \dataMemory[31][14] ;
 wire \dataMemory[31][15] ;
 wire \dataMemory[31][16] ;
 wire \dataMemory[31][17] ;
 wire \dataMemory[31][18] ;
 wire \dataMemory[31][19] ;
 wire \dataMemory[31][1] ;
 wire \dataMemory[31][20] ;
 wire \dataMemory[31][21] ;
 wire \dataMemory[31][22] ;
 wire \dataMemory[31][23] ;
 wire \dataMemory[31][24] ;
 wire \dataMemory[31][25] ;
 wire \dataMemory[31][26] ;
 wire \dataMemory[31][27] ;
 wire \dataMemory[31][28] ;
 wire \dataMemory[31][29] ;
 wire \dataMemory[31][2] ;
 wire \dataMemory[31][30] ;
 wire \dataMemory[31][31] ;
 wire \dataMemory[31][3] ;
 wire \dataMemory[31][4] ;
 wire \dataMemory[31][5] ;
 wire \dataMemory[31][6] ;
 wire \dataMemory[31][7] ;
 wire \dataMemory[31][8] ;
 wire \dataMemory[31][9] ;
 wire \dataMemory[3][0] ;
 wire \dataMemory[3][10] ;
 wire \dataMemory[3][11] ;
 wire \dataMemory[3][12] ;
 wire \dataMemory[3][13] ;
 wire \dataMemory[3][14] ;
 wire \dataMemory[3][15] ;
 wire \dataMemory[3][16] ;
 wire \dataMemory[3][17] ;
 wire \dataMemory[3][18] ;
 wire \dataMemory[3][19] ;
 wire \dataMemory[3][1] ;
 wire \dataMemory[3][20] ;
 wire \dataMemory[3][21] ;
 wire \dataMemory[3][22] ;
 wire \dataMemory[3][23] ;
 wire \dataMemory[3][24] ;
 wire \dataMemory[3][25] ;
 wire \dataMemory[3][26] ;
 wire \dataMemory[3][27] ;
 wire \dataMemory[3][28] ;
 wire \dataMemory[3][29] ;
 wire \dataMemory[3][2] ;
 wire \dataMemory[3][30] ;
 wire \dataMemory[3][31] ;
 wire \dataMemory[3][3] ;
 wire \dataMemory[3][4] ;
 wire \dataMemory[3][5] ;
 wire \dataMemory[3][6] ;
 wire \dataMemory[3][7] ;
 wire \dataMemory[3][8] ;
 wire \dataMemory[3][9] ;
 wire \dataMemory[4][0] ;
 wire \dataMemory[4][10] ;
 wire \dataMemory[4][11] ;
 wire \dataMemory[4][12] ;
 wire \dataMemory[4][13] ;
 wire \dataMemory[4][14] ;
 wire \dataMemory[4][15] ;
 wire \dataMemory[4][16] ;
 wire \dataMemory[4][17] ;
 wire \dataMemory[4][18] ;
 wire \dataMemory[4][19] ;
 wire \dataMemory[4][1] ;
 wire \dataMemory[4][20] ;
 wire \dataMemory[4][21] ;
 wire \dataMemory[4][22] ;
 wire \dataMemory[4][23] ;
 wire \dataMemory[4][24] ;
 wire \dataMemory[4][25] ;
 wire \dataMemory[4][26] ;
 wire \dataMemory[4][27] ;
 wire \dataMemory[4][28] ;
 wire \dataMemory[4][29] ;
 wire \dataMemory[4][2] ;
 wire \dataMemory[4][30] ;
 wire \dataMemory[4][31] ;
 wire \dataMemory[4][3] ;
 wire \dataMemory[4][4] ;
 wire \dataMemory[4][5] ;
 wire \dataMemory[4][6] ;
 wire \dataMemory[4][7] ;
 wire \dataMemory[4][8] ;
 wire \dataMemory[4][9] ;
 wire \dataMemory[5][0] ;
 wire \dataMemory[5][10] ;
 wire \dataMemory[5][11] ;
 wire \dataMemory[5][12] ;
 wire \dataMemory[5][13] ;
 wire \dataMemory[5][14] ;
 wire \dataMemory[5][15] ;
 wire \dataMemory[5][16] ;
 wire \dataMemory[5][17] ;
 wire \dataMemory[5][18] ;
 wire \dataMemory[5][19] ;
 wire \dataMemory[5][1] ;
 wire \dataMemory[5][20] ;
 wire \dataMemory[5][21] ;
 wire \dataMemory[5][22] ;
 wire \dataMemory[5][23] ;
 wire \dataMemory[5][24] ;
 wire \dataMemory[5][25] ;
 wire \dataMemory[5][26] ;
 wire \dataMemory[5][27] ;
 wire \dataMemory[5][28] ;
 wire \dataMemory[5][29] ;
 wire \dataMemory[5][2] ;
 wire \dataMemory[5][30] ;
 wire \dataMemory[5][31] ;
 wire \dataMemory[5][3] ;
 wire \dataMemory[5][4] ;
 wire \dataMemory[5][5] ;
 wire \dataMemory[5][6] ;
 wire \dataMemory[5][7] ;
 wire \dataMemory[5][8] ;
 wire \dataMemory[5][9] ;
 wire \dataMemory[6][0] ;
 wire \dataMemory[6][10] ;
 wire \dataMemory[6][11] ;
 wire \dataMemory[6][12] ;
 wire \dataMemory[6][13] ;
 wire \dataMemory[6][14] ;
 wire \dataMemory[6][15] ;
 wire \dataMemory[6][16] ;
 wire \dataMemory[6][17] ;
 wire \dataMemory[6][18] ;
 wire \dataMemory[6][19] ;
 wire \dataMemory[6][1] ;
 wire \dataMemory[6][20] ;
 wire \dataMemory[6][21] ;
 wire \dataMemory[6][22] ;
 wire \dataMemory[6][23] ;
 wire \dataMemory[6][24] ;
 wire \dataMemory[6][25] ;
 wire \dataMemory[6][26] ;
 wire \dataMemory[6][27] ;
 wire \dataMemory[6][28] ;
 wire \dataMemory[6][29] ;
 wire \dataMemory[6][2] ;
 wire \dataMemory[6][30] ;
 wire \dataMemory[6][31] ;
 wire \dataMemory[6][3] ;
 wire \dataMemory[6][4] ;
 wire \dataMemory[6][5] ;
 wire \dataMemory[6][6] ;
 wire \dataMemory[6][7] ;
 wire \dataMemory[6][8] ;
 wire \dataMemory[6][9] ;
 wire \dataMemory[7][0] ;
 wire \dataMemory[7][10] ;
 wire \dataMemory[7][11] ;
 wire \dataMemory[7][12] ;
 wire \dataMemory[7][13] ;
 wire \dataMemory[7][14] ;
 wire \dataMemory[7][15] ;
 wire \dataMemory[7][16] ;
 wire \dataMemory[7][17] ;
 wire \dataMemory[7][18] ;
 wire \dataMemory[7][19] ;
 wire \dataMemory[7][1] ;
 wire \dataMemory[7][20] ;
 wire \dataMemory[7][21] ;
 wire \dataMemory[7][22] ;
 wire \dataMemory[7][23] ;
 wire \dataMemory[7][24] ;
 wire \dataMemory[7][25] ;
 wire \dataMemory[7][26] ;
 wire \dataMemory[7][27] ;
 wire \dataMemory[7][28] ;
 wire \dataMemory[7][29] ;
 wire \dataMemory[7][2] ;
 wire \dataMemory[7][30] ;
 wire \dataMemory[7][31] ;
 wire \dataMemory[7][3] ;
 wire \dataMemory[7][4] ;
 wire \dataMemory[7][5] ;
 wire \dataMemory[7][6] ;
 wire \dataMemory[7][7] ;
 wire \dataMemory[7][8] ;
 wire \dataMemory[7][9] ;
 wire \dataMemory[8][0] ;
 wire \dataMemory[8][10] ;
 wire \dataMemory[8][11] ;
 wire \dataMemory[8][12] ;
 wire \dataMemory[8][13] ;
 wire \dataMemory[8][14] ;
 wire \dataMemory[8][15] ;
 wire \dataMemory[8][16] ;
 wire \dataMemory[8][17] ;
 wire \dataMemory[8][18] ;
 wire \dataMemory[8][19] ;
 wire \dataMemory[8][1] ;
 wire \dataMemory[8][20] ;
 wire \dataMemory[8][21] ;
 wire \dataMemory[8][22] ;
 wire \dataMemory[8][23] ;
 wire \dataMemory[8][24] ;
 wire \dataMemory[8][25] ;
 wire \dataMemory[8][26] ;
 wire \dataMemory[8][27] ;
 wire \dataMemory[8][28] ;
 wire \dataMemory[8][29] ;
 wire \dataMemory[8][2] ;
 wire \dataMemory[8][30] ;
 wire \dataMemory[8][31] ;
 wire \dataMemory[8][3] ;
 wire \dataMemory[8][4] ;
 wire \dataMemory[8][5] ;
 wire \dataMemory[8][6] ;
 wire \dataMemory[8][7] ;
 wire \dataMemory[8][8] ;
 wire \dataMemory[8][9] ;
 wire \dataMemory[9][0] ;
 wire \dataMemory[9][10] ;
 wire \dataMemory[9][11] ;
 wire \dataMemory[9][12] ;
 wire \dataMemory[9][13] ;
 wire \dataMemory[9][14] ;
 wire \dataMemory[9][15] ;
 wire \dataMemory[9][16] ;
 wire \dataMemory[9][17] ;
 wire \dataMemory[9][18] ;
 wire \dataMemory[9][19] ;
 wire \dataMemory[9][1] ;
 wire \dataMemory[9][20] ;
 wire \dataMemory[9][21] ;
 wire \dataMemory[9][22] ;
 wire \dataMemory[9][23] ;
 wire \dataMemory[9][24] ;
 wire \dataMemory[9][25] ;
 wire \dataMemory[9][26] ;
 wire \dataMemory[9][27] ;
 wire \dataMemory[9][28] ;
 wire \dataMemory[9][29] ;
 wire \dataMemory[9][2] ;
 wire \dataMemory[9][30] ;
 wire \dataMemory[9][31] ;
 wire \dataMemory[9][3] ;
 wire \dataMemory[9][4] ;
 wire \dataMemory[9][5] ;
 wire \dataMemory[9][6] ;
 wire \dataMemory[9][7] ;
 wire \dataMemory[9][8] ;
 wire \dataMemory[9][9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__1845__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A_N (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__B (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__S0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__C (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__S0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__S1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__S0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__S0 (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__S0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__S1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__S0 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__S1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__C1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__C1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__S1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__S1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S0 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__S1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2001__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__S1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__S0 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__S1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2031__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2031__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__S0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__S1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__S0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__S1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__S0 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__S1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__B (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__C1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__S1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2079__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2079__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__S0 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__S1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__S1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__S1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__S0 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__S1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__S0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__S1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__S1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__S1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__S1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__C1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__S0 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__S1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__A1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__S0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__S1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__B (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__S0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__S1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__S0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__S1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__S0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__S1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__A1 (.DIODE(_1438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__S0 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__S1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__S0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__S1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__S0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__S1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__S1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__S0 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__S1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__S1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__S (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__S0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__S1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__S0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__S1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__S0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__S1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__S0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__S1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S0 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__C1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__C1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__S0 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__S1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__S0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__S1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__S0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__S1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__S0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__S1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__S0 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__S1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__S0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__S1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__B (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__B (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__C1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__S0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__S1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__S1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__S1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__S0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__S1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__C1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__S0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__S1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A1 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__S0 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__S1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__S0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__S1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__S (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__B (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__C1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__S1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__C1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__B (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__C1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__S0 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__S1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A_N (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__C (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__B (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__A0 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__S (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__S (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__C_N (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2714__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__S (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__S (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__S (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__S (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__S (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__C (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2854__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2863__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2866__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__S (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2883__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2894__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2904__S (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2917__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2917__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__A0 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2930__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__S (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__S (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__C (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A0 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__S (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__S (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__S (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__S (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__S (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__S (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__S (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__S (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__C (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__S (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__S (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__S (.DIODE(_1831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__S (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__S (.DIODE(_1833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__S (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__S (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__S (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__S (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A0 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A0 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A0 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A0 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__S (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__S (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__S (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__S (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__S (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__S (.DIODE(_1840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__S (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__S (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__S (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__S (.DIODE(_1842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__S (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__S (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__S (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__S (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A0 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A0 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A0 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__S (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__S (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__CLK (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__CLK (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__CLK (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__CLK (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__CLK (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__CLK (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__CLK (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__CLK (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__CLK (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__CLK (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__CLK (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__CLK (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__CLK (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__CLK (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__CLK (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__CLK (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__CLK (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__CLK (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__CLK (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__CLK (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__CLK (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__CLK (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__CLK (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__CLK (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__CLK (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__CLK (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__CLK (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__CLK (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__CLK (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__CLK (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__CLK (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__CLK (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_1813_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(_1813_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(_1812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(_1838_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_1835_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout339_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout362_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout378_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout380_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout387_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net389));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(_1842_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(_1840_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_1839_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_1833_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_1832_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(_1831_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_980 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_998 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _1845_ (.A(net212),
    .Y(_1024_));
 sky130_fd_sc_hd__inv_4 _1846_ (.A(net206),
    .Y(_1025_));
 sky130_fd_sc_hd__nor2_1 _1847_ (.A(net280),
    .B(net242),
    .Y(_1026_));
 sky130_fd_sc_hd__and2b_1 _1848_ (.A_N(net281),
    .B(net243),
    .X(_1027_));
 sky130_fd_sc_hd__and2b_1 _1849_ (.A_N(net242),
    .B(net280),
    .X(_1028_));
 sky130_fd_sc_hd__and3_1 _1850_ (.A(net278),
    .B(net240),
    .C(\dataMemory[23][0] ),
    .X(_1029_));
 sky130_fd_sc_hd__a221o_1 _1851_ (.A1(\dataMemory[22][0] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[21][0] ),
    .C1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__a211o_1 _1852_ (.A1(\dataMemory[20][0] ),
    .A2(net167),
    .B1(_1030_),
    .C1(net187),
    .X(_1031_));
 sky130_fd_sc_hd__and3_1 _1853_ (.A(net278),
    .B(net240),
    .C(\dataMemory[19][0] ),
    .X(_1032_));
 sky130_fd_sc_hd__a221o_1 _1854_ (.A1(\dataMemory[18][0] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[17][0] ),
    .C1(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__a211o_1 _1855_ (.A1(\dataMemory[16][0] ),
    .A2(net167),
    .B1(_1033_),
    .C1(net211),
    .X(_1034_));
 sky130_fd_sc_hd__and3_1 _1856_ (.A(net278),
    .B(net240),
    .C(\dataMemory[27][0] ),
    .X(_1035_));
 sky130_fd_sc_hd__a221o_1 _1857_ (.A1(\dataMemory[24][0] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[25][0] ),
    .C1(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__a211o_1 _1858_ (.A1(\dataMemory[26][0] ),
    .A2(net151),
    .B1(_1036_),
    .C1(net211),
    .X(_1037_));
 sky130_fd_sc_hd__mux4_1 _1859_ (.A0(\dataMemory[28][0] ),
    .A1(\dataMemory[29][0] ),
    .A2(\dataMemory[30][0] ),
    .A3(\dataMemory[31][0] ),
    .S0(net278),
    .S1(net240),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_2 _1860_ (.A(net208),
    .B(net204),
    .Y(_1039_));
 sky130_fd_sc_hd__and3_1 _1861_ (.A(net279),
    .B(net241),
    .C(\dataMemory[7][0] ),
    .X(_1040_));
 sky130_fd_sc_hd__a221o_1 _1862_ (.A1(\dataMemory[6][0] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[5][0] ),
    .C1(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__a211o_1 _1863_ (.A1(\dataMemory[4][0] ),
    .A2(net168),
    .B1(_1041_),
    .C1(net196),
    .X(_1042_));
 sky130_fd_sc_hd__and3_1 _1864_ (.A(net279),
    .B(\dataMemory[3][0] ),
    .C(net241),
    .X(_1043_));
 sky130_fd_sc_hd__a221o_1 _1865_ (.A1(\dataMemory[2][0] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[1][0] ),
    .C1(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__a211o_1 _1866_ (.A1(\dataMemory[0][0] ),
    .A2(net168),
    .B1(_1044_),
    .C1(net211),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _1867_ (.A(net208),
    .B(net204),
    .Y(_1046_));
 sky130_fd_sc_hd__and3_1 _1868_ (.A(net278),
    .B(net240),
    .C(\dataMemory[11][0] ),
    .X(_1047_));
 sky130_fd_sc_hd__a221o_1 _1869_ (.A1(\dataMemory[8][0] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[9][0] ),
    .C1(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__a211o_1 _1870_ (.A1(\dataMemory[10][0] ),
    .A2(net152),
    .B1(_1048_),
    .C1(net211),
    .X(_1049_));
 sky130_fd_sc_hd__mux4_1 _1871_ (.A0(\dataMemory[12][0] ),
    .A1(\dataMemory[13][0] ),
    .A2(\dataMemory[14][0] ),
    .A3(\dataMemory[15][0] ),
    .S0(net279),
    .S1(net241),
    .X(_1050_));
 sky130_fd_sc_hd__o21a_1 _1872_ (.A1(net187),
    .A2(_1050_),
    .B1(net206),
    .X(_1051_));
 sky130_fd_sc_hd__a32o_1 _1873_ (.A1(net183),
    .A2(_1042_),
    .A3(_1045_),
    .B1(_1049_),
    .B2(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__o21a_1 _1874_ (.A1(net187),
    .A2(_1038_),
    .B1(net206),
    .X(_1053_));
 sky130_fd_sc_hd__a32o_1 _1875_ (.A1(net183),
    .A2(_1031_),
    .A3(_1034_),
    .B1(_1037_),
    .B2(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__mux2_4 _1876_ (.A0(_1052_),
    .A1(_1054_),
    .S(net203),
    .X(net40));
 sky130_fd_sc_hd__and3_1 _1877_ (.A(net278),
    .B(net240),
    .C(\dataMemory[23][1] ),
    .X(_1055_));
 sky130_fd_sc_hd__a221o_1 _1878_ (.A1(\dataMemory[22][1] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[21][1] ),
    .C1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__a211o_1 _1879_ (.A1(\dataMemory[20][1] ),
    .A2(net167),
    .B1(_1056_),
    .C1(net187),
    .X(_1057_));
 sky130_fd_sc_hd__and3_1 _1880_ (.A(net278),
    .B(net240),
    .C(\dataMemory[19][1] ),
    .X(_1058_));
 sky130_fd_sc_hd__a221o_1 _1881_ (.A1(\dataMemory[18][1] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[17][1] ),
    .C1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__a211o_1 _1882_ (.A1(\dataMemory[16][1] ),
    .A2(net167),
    .B1(_1059_),
    .C1(net211),
    .X(_1060_));
 sky130_fd_sc_hd__and3_1 _1883_ (.A(net278),
    .B(net240),
    .C(\dataMemory[27][1] ),
    .X(_1061_));
 sky130_fd_sc_hd__a221o_1 _1884_ (.A1(\dataMemory[24][1] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[25][1] ),
    .C1(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__a211o_1 _1885_ (.A1(\dataMemory[26][1] ),
    .A2(net151),
    .B1(_1062_),
    .C1(net211),
    .X(_1063_));
 sky130_fd_sc_hd__mux4_1 _1886_ (.A0(\dataMemory[28][1] ),
    .A1(\dataMemory[29][1] ),
    .A2(\dataMemory[30][1] ),
    .A3(\dataMemory[31][1] ),
    .S0(net278),
    .S1(net240),
    .X(_1064_));
 sky130_fd_sc_hd__and3_1 _1887_ (.A(net279),
    .B(net241),
    .C(\dataMemory[7][1] ),
    .X(_1065_));
 sky130_fd_sc_hd__a221o_1 _1888_ (.A1(\dataMemory[6][1] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[5][1] ),
    .C1(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__a211o_1 _1889_ (.A1(\dataMemory[4][1] ),
    .A2(net168),
    .B1(_1066_),
    .C1(net187),
    .X(_1067_));
 sky130_fd_sc_hd__and3_1 _1890_ (.A(net279),
    .B(net241),
    .C(\dataMemory[3][1] ),
    .X(_1068_));
 sky130_fd_sc_hd__a221o_1 _1891_ (.A1(\dataMemory[2][1] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[1][1] ),
    .C1(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__a211o_1 _1892_ (.A1(\dataMemory[0][1] ),
    .A2(net168),
    .B1(_1069_),
    .C1(net211),
    .X(_1070_));
 sky130_fd_sc_hd__and3_1 _1893_ (.A(net279),
    .B(net241),
    .C(\dataMemory[11][1] ),
    .X(_1071_));
 sky130_fd_sc_hd__a221o_1 _1894_ (.A1(\dataMemory[8][1] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[9][1] ),
    .C1(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__a211o_1 _1895_ (.A1(\dataMemory[10][1] ),
    .A2(net151),
    .B1(_1072_),
    .C1(net211),
    .X(_1073_));
 sky130_fd_sc_hd__mux4_1 _1896_ (.A0(\dataMemory[12][1] ),
    .A1(\dataMemory[13][1] ),
    .A2(\dataMemory[14][1] ),
    .A3(\dataMemory[15][1] ),
    .S0(net279),
    .S1(net241),
    .X(_1074_));
 sky130_fd_sc_hd__o21a_1 _1897_ (.A1(net187),
    .A2(_1074_),
    .B1(net206),
    .X(_1075_));
 sky130_fd_sc_hd__a32o_1 _1898_ (.A1(net183),
    .A2(_1067_),
    .A3(_1070_),
    .B1(_1073_),
    .B2(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__o21a_1 _1899_ (.A1(net187),
    .A2(_1064_),
    .B1(net206),
    .X(_1077_));
 sky130_fd_sc_hd__a32o_1 _1900_ (.A1(net183),
    .A2(_1057_),
    .A3(_1060_),
    .B1(_1063_),
    .B2(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_4 _1901_ (.A0(_1076_),
    .A1(_1078_),
    .S(net203),
    .X(net51));
 sky130_fd_sc_hd__and3_1 _1902_ (.A(net278),
    .B(net240),
    .C(\dataMemory[23][2] ),
    .X(_1079_));
 sky130_fd_sc_hd__a221o_1 _1903_ (.A1(\dataMemory[22][2] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[21][2] ),
    .C1(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__a211o_1 _1904_ (.A1(\dataMemory[20][2] ),
    .A2(net167),
    .B1(_1080_),
    .C1(net187),
    .X(_1081_));
 sky130_fd_sc_hd__and3_1 _1905_ (.A(net278),
    .B(net240),
    .C(\dataMemory[19][2] ),
    .X(_1082_));
 sky130_fd_sc_hd__a221o_1 _1906_ (.A1(\dataMemory[18][2] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[17][2] ),
    .C1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__a211o_1 _1907_ (.A1(\dataMemory[16][2] ),
    .A2(net167),
    .B1(_1083_),
    .C1(net211),
    .X(_1084_));
 sky130_fd_sc_hd__and3_1 _1908_ (.A(net278),
    .B(net240),
    .C(\dataMemory[27][2] ),
    .X(_1085_));
 sky130_fd_sc_hd__a221o_1 _1909_ (.A1(\dataMemory[24][2] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[25][2] ),
    .C1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__a211o_1 _1910_ (.A1(\dataMemory[26][2] ),
    .A2(net151),
    .B1(_1086_),
    .C1(net211),
    .X(_1087_));
 sky130_fd_sc_hd__mux4_1 _1911_ (.A0(\dataMemory[28][2] ),
    .A1(\dataMemory[29][2] ),
    .A2(\dataMemory[30][2] ),
    .A3(\dataMemory[31][2] ),
    .S0(net278),
    .S1(net240),
    .X(_1088_));
 sky130_fd_sc_hd__and3_1 _1912_ (.A(net279),
    .B(net241),
    .C(\dataMemory[7][2] ),
    .X(_1089_));
 sky130_fd_sc_hd__a221o_1 _1913_ (.A1(\dataMemory[6][2] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[5][2] ),
    .C1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__a211o_1 _1914_ (.A1(\dataMemory[4][2] ),
    .A2(net168),
    .B1(_1090_),
    .C1(net187),
    .X(_1091_));
 sky130_fd_sc_hd__and3_1 _1915_ (.A(net279),
    .B(net241),
    .C(\dataMemory[3][2] ),
    .X(_1092_));
 sky130_fd_sc_hd__a221o_1 _1916_ (.A1(\dataMemory[2][2] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[1][2] ),
    .C1(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__a211o_1 _1917_ (.A1(\dataMemory[0][2] ),
    .A2(net168),
    .B1(_1093_),
    .C1(net211),
    .X(_1094_));
 sky130_fd_sc_hd__and3_1 _1918_ (.A(net279),
    .B(net241),
    .C(\dataMemory[11][2] ),
    .X(_1095_));
 sky130_fd_sc_hd__a221o_1 _1919_ (.A1(\dataMemory[8][2] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[9][2] ),
    .C1(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__a211o_1 _1920_ (.A1(\dataMemory[10][2] ),
    .A2(net151),
    .B1(_1096_),
    .C1(net211),
    .X(_1097_));
 sky130_fd_sc_hd__mux4_1 _1921_ (.A0(\dataMemory[12][2] ),
    .A1(\dataMemory[13][2] ),
    .A2(\dataMemory[14][2] ),
    .A3(\dataMemory[15][2] ),
    .S0(net279),
    .S1(net241),
    .X(_1098_));
 sky130_fd_sc_hd__o21a_1 _1922_ (.A1(net187),
    .A2(_1098_),
    .B1(net206),
    .X(_1099_));
 sky130_fd_sc_hd__a32o_1 _1923_ (.A1(net183),
    .A2(_1091_),
    .A3(_1094_),
    .B1(_1097_),
    .B2(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__o21a_1 _1924_ (.A1(net187),
    .A2(_1088_),
    .B1(net206),
    .X(_1101_));
 sky130_fd_sc_hd__a32o_1 _1925_ (.A1(net183),
    .A2(_1081_),
    .A3(_1084_),
    .B1(_1087_),
    .B2(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__mux2_4 _1926_ (.A0(_1100_),
    .A1(_1102_),
    .S(net203),
    .X(net62));
 sky130_fd_sc_hd__and3_1 _1927_ (.A(net278),
    .B(net240),
    .C(\dataMemory[23][3] ),
    .X(_1103_));
 sky130_fd_sc_hd__a221o_1 _1928_ (.A1(\dataMemory[22][3] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[21][3] ),
    .C1(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__a211o_1 _1929_ (.A1(\dataMemory[20][3] ),
    .A2(net167),
    .B1(_1104_),
    .C1(net187),
    .X(_1105_));
 sky130_fd_sc_hd__and3_1 _1930_ (.A(net278),
    .B(net240),
    .C(\dataMemory[19][3] ),
    .X(_1106_));
 sky130_fd_sc_hd__a221o_1 _1931_ (.A1(\dataMemory[18][3] ),
    .A2(net151),
    .B1(net136),
    .B2(\dataMemory[17][3] ),
    .C1(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__a211o_1 _1932_ (.A1(\dataMemory[16][3] ),
    .A2(net167),
    .B1(_1107_),
    .C1(net211),
    .X(_1108_));
 sky130_fd_sc_hd__and3_1 _1933_ (.A(net278),
    .B(net240),
    .C(\dataMemory[27][3] ),
    .X(_1109_));
 sky130_fd_sc_hd__a221o_1 _1934_ (.A1(\dataMemory[24][3] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[25][3] ),
    .C1(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a211o_1 _1935_ (.A1(\dataMemory[26][3] ),
    .A2(net151),
    .B1(_1110_),
    .C1(net211),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_1 _1936_ (.A0(\dataMemory[28][3] ),
    .A1(\dataMemory[29][3] ),
    .A2(\dataMemory[30][3] ),
    .A3(\dataMemory[31][3] ),
    .S0(net279),
    .S1(net248),
    .X(_1112_));
 sky130_fd_sc_hd__and3_1 _1937_ (.A(net279),
    .B(net241),
    .C(\dataMemory[7][3] ),
    .X(_1113_));
 sky130_fd_sc_hd__a221o_1 _1938_ (.A1(\dataMemory[6][3] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[5][3] ),
    .C1(_1113_),
    .X(_1114_));
 sky130_fd_sc_hd__a211o_1 _1939_ (.A1(\dataMemory[4][3] ),
    .A2(net168),
    .B1(_1114_),
    .C1(net187),
    .X(_1115_));
 sky130_fd_sc_hd__and3_1 _1940_ (.A(net279),
    .B(net241),
    .C(\dataMemory[3][3] ),
    .X(_1116_));
 sky130_fd_sc_hd__a221o_1 _1941_ (.A1(\dataMemory[2][3] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[1][3] ),
    .C1(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__a211o_1 _1942_ (.A1(\dataMemory[0][3] ),
    .A2(net168),
    .B1(_1117_),
    .C1(net211),
    .X(_1118_));
 sky130_fd_sc_hd__and3_1 _1943_ (.A(net279),
    .B(net241),
    .C(\dataMemory[11][3] ),
    .X(_1119_));
 sky130_fd_sc_hd__a221o_1 _1944_ (.A1(\dataMemory[8][3] ),
    .A2(net167),
    .B1(net136),
    .B2(\dataMemory[9][3] ),
    .C1(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__a211o_1 _1945_ (.A1(\dataMemory[10][3] ),
    .A2(net151),
    .B1(_1120_),
    .C1(net211),
    .X(_1121_));
 sky130_fd_sc_hd__mux4_1 _1946_ (.A0(\dataMemory[12][3] ),
    .A1(\dataMemory[13][3] ),
    .A2(\dataMemory[14][3] ),
    .A3(\dataMemory[15][3] ),
    .S0(net286),
    .S1(net241),
    .X(_1122_));
 sky130_fd_sc_hd__o21a_1 _1947_ (.A1(net187),
    .A2(_1122_),
    .B1(net206),
    .X(_1123_));
 sky130_fd_sc_hd__a32o_1 _1948_ (.A1(net183),
    .A2(_1115_),
    .A3(_1118_),
    .B1(_1121_),
    .B2(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__o21a_1 _1949_ (.A1(net187),
    .A2(_1112_),
    .B1(net206),
    .X(_1125_));
 sky130_fd_sc_hd__a32o_1 _1950_ (.A1(net183),
    .A2(_1105_),
    .A3(_1108_),
    .B1(_1111_),
    .B2(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_4 _1951_ (.A0(_1124_),
    .A1(_1126_),
    .S(net203),
    .X(net65));
 sky130_fd_sc_hd__and3_1 _1952_ (.A(net282),
    .B(net244),
    .C(\dataMemory[23][4] ),
    .X(_1127_));
 sky130_fd_sc_hd__a221o_1 _1953_ (.A1(\dataMemory[22][4] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[21][4] ),
    .C1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__a211o_1 _1954_ (.A1(\dataMemory[20][4] ),
    .A2(net171),
    .B1(_1128_),
    .C1(net189),
    .X(_1129_));
 sky130_fd_sc_hd__and3_1 _1955_ (.A(net282),
    .B(net244),
    .C(\dataMemory[19][4] ),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_1 _1956_ (.A1(\dataMemory[18][4] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[17][4] ),
    .C1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__a211o_1 _1957_ (.A1(\dataMemory[16][4] ),
    .A2(net171),
    .B1(_1131_),
    .C1(net213),
    .X(_1132_));
 sky130_fd_sc_hd__and3_1 _1958_ (.A(net286),
    .B(net241),
    .C(\dataMemory[27][4] ),
    .X(_1133_));
 sky130_fd_sc_hd__a221o_1 _1959_ (.A1(\dataMemory[24][4] ),
    .A2(net168),
    .B1(net137),
    .B2(\dataMemory[25][4] ),
    .C1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__a211o_1 _1960_ (.A1(\dataMemory[26][4] ),
    .A2(net152),
    .B1(_1134_),
    .C1(net215),
    .X(_1135_));
 sky130_fd_sc_hd__mux4_1 _1961_ (.A0(\dataMemory[28][4] ),
    .A1(\dataMemory[29][4] ),
    .A2(\dataMemory[30][4] ),
    .A3(\dataMemory[31][4] ),
    .S0(net282),
    .S1(net244),
    .X(_1136_));
 sky130_fd_sc_hd__and3_1 _1962_ (.A(net282),
    .B(net244),
    .C(\dataMemory[7][4] ),
    .X(_1137_));
 sky130_fd_sc_hd__a221o_1 _1963_ (.A1(\dataMemory[6][4] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[5][4] ),
    .C1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__a211o_1 _1964_ (.A1(\dataMemory[4][4] ),
    .A2(net171),
    .B1(_1138_),
    .C1(net189),
    .X(_1139_));
 sky130_fd_sc_hd__and3_1 _1965_ (.A(net282),
    .B(net244),
    .C(\dataMemory[3][4] ),
    .X(_1140_));
 sky130_fd_sc_hd__a221o_1 _1966_ (.A1(\dataMemory[2][4] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[1][4] ),
    .C1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__a211o_1 _1967_ (.A1(\dataMemory[0][4] ),
    .A2(net171),
    .B1(_1141_),
    .C1(net213),
    .X(_1142_));
 sky130_fd_sc_hd__and3_1 _1968_ (.A(net282),
    .B(net244),
    .C(\dataMemory[11][4] ),
    .X(_1143_));
 sky130_fd_sc_hd__a221o_1 _1969_ (.A1(\dataMemory[8][4] ),
    .A2(net168),
    .B1(net137),
    .B2(\dataMemory[9][4] ),
    .C1(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__a211o_1 _1970_ (.A1(\dataMemory[10][4] ),
    .A2(net151),
    .B1(_1144_),
    .C1(net215),
    .X(_1145_));
 sky130_fd_sc_hd__mux4_1 _1971_ (.A0(\dataMemory[12][4] ),
    .A1(\dataMemory[13][4] ),
    .A2(\dataMemory[14][4] ),
    .A3(\dataMemory[15][4] ),
    .S0(net282),
    .S1(net244),
    .X(_1146_));
 sky130_fd_sc_hd__o21a_1 _1972_ (.A1(net189),
    .A2(_1146_),
    .B1(net207),
    .X(_1147_));
 sky130_fd_sc_hd__a32o_1 _1973_ (.A1(net184),
    .A2(_1139_),
    .A3(_1142_),
    .B1(_1145_),
    .B2(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__o21a_1 _1974_ (.A1(net187),
    .A2(_1136_),
    .B1(net207),
    .X(_1149_));
 sky130_fd_sc_hd__a32o_1 _1975_ (.A1(net184),
    .A2(_1129_),
    .A3(_1132_),
    .B1(_1135_),
    .B2(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_4 _1976_ (.A0(_1148_),
    .A1(_1150_),
    .S(net203),
    .X(net66));
 sky130_fd_sc_hd__and3_1 _1977_ (.A(net280),
    .B(net242),
    .C(\dataMemory[23][5] ),
    .X(_1151_));
 sky130_fd_sc_hd__a221o_1 _1978_ (.A1(\dataMemory[22][5] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[21][5] ),
    .C1(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__a211o_1 _1979_ (.A1(\dataMemory[20][5] ),
    .A2(net169),
    .B1(_1152_),
    .C1(net188),
    .X(_1153_));
 sky130_fd_sc_hd__and3_1 _1980_ (.A(net280),
    .B(net242),
    .C(\dataMemory[19][5] ),
    .X(_1154_));
 sky130_fd_sc_hd__a221o_1 _1981_ (.A1(\dataMemory[18][5] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[17][5] ),
    .C1(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__a211o_1 _1982_ (.A1(\dataMemory[16][5] ),
    .A2(net169),
    .B1(_1155_),
    .C1(net212),
    .X(_1156_));
 sky130_fd_sc_hd__and3_1 _1983_ (.A(net280),
    .B(net242),
    .C(\dataMemory[27][5] ),
    .X(_1157_));
 sky130_fd_sc_hd__a221o_1 _1984_ (.A1(\dataMemory[24][5] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[25][5] ),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__a211o_1 _1985_ (.A1(\dataMemory[26][5] ),
    .A2(net153),
    .B1(_1158_),
    .C1(net212),
    .X(_1159_));
 sky130_fd_sc_hd__mux4_1 _1986_ (.A0(\dataMemory[28][5] ),
    .A1(\dataMemory[29][5] ),
    .A2(\dataMemory[30][5] ),
    .A3(\dataMemory[31][5] ),
    .S0(net280),
    .S1(net242),
    .X(_1160_));
 sky130_fd_sc_hd__and3_1 _1987_ (.A(net281),
    .B(net243),
    .C(\dataMemory[7][5] ),
    .X(_1161_));
 sky130_fd_sc_hd__a221o_1 _1988_ (.A1(\dataMemory[6][5] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[5][5] ),
    .C1(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__a211o_1 _1989_ (.A1(\dataMemory[4][5] ),
    .A2(net170),
    .B1(_1162_),
    .C1(net188),
    .X(_1163_));
 sky130_fd_sc_hd__and3_1 _1990_ (.A(net281),
    .B(net243),
    .C(\dataMemory[3][5] ),
    .X(_1164_));
 sky130_fd_sc_hd__a221o_1 _1991_ (.A1(\dataMemory[2][5] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[1][5] ),
    .C1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__a211o_1 _1992_ (.A1(\dataMemory[0][5] ),
    .A2(net170),
    .B1(_1165_),
    .C1(net212),
    .X(_1166_));
 sky130_fd_sc_hd__and3_1 _1993_ (.A(net280),
    .B(net242),
    .C(\dataMemory[11][5] ),
    .X(_1167_));
 sky130_fd_sc_hd__a221o_1 _1994_ (.A1(\dataMemory[8][5] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[9][5] ),
    .C1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__a211o_1 _1995_ (.A1(\dataMemory[10][5] ),
    .A2(net153),
    .B1(_1168_),
    .C1(net212),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_1 _1996_ (.A0(\dataMemory[12][5] ),
    .A1(\dataMemory[13][5] ),
    .A2(\dataMemory[14][5] ),
    .A3(\dataMemory[15][5] ),
    .S0(net281),
    .S1(net243),
    .X(_1170_));
 sky130_fd_sc_hd__o21a_1 _1997_ (.A1(net188),
    .A2(_1170_),
    .B1(net206),
    .X(_1171_));
 sky130_fd_sc_hd__a32o_1 _1998_ (.A1(net183),
    .A2(_1163_),
    .A3(_1166_),
    .B1(_1169_),
    .B2(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__o21a_1 _1999_ (.A1(net188),
    .A2(_1160_),
    .B1(net206),
    .X(_1173_));
 sky130_fd_sc_hd__a32o_1 _2000_ (.A1(net184),
    .A2(_1153_),
    .A3(_1156_),
    .B1(_1159_),
    .B2(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__mux2_4 _2001_ (.A0(_1172_),
    .A1(_1174_),
    .S(net203),
    .X(net67));
 sky130_fd_sc_hd__and3_1 _2002_ (.A(net282),
    .B(net244),
    .C(\dataMemory[23][6] ),
    .X(_1175_));
 sky130_fd_sc_hd__a221o_1 _2003_ (.A1(\dataMemory[22][6] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[21][6] ),
    .C1(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__a211o_1 _2004_ (.A1(\dataMemory[20][6] ),
    .A2(net171),
    .B1(_1176_),
    .C1(net189),
    .X(_1177_));
 sky130_fd_sc_hd__and3_1 _2005_ (.A(net282),
    .B(net244),
    .C(\dataMemory[19][6] ),
    .X(_1178_));
 sky130_fd_sc_hd__a221o_1 _2006_ (.A1(\dataMemory[18][6] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[17][6] ),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__a211o_1 _2007_ (.A1(\dataMemory[16][6] ),
    .A2(net171),
    .B1(_1179_),
    .C1(net213),
    .X(_1180_));
 sky130_fd_sc_hd__and3_1 _2008_ (.A(net282),
    .B(net244),
    .C(\dataMemory[27][6] ),
    .X(_1181_));
 sky130_fd_sc_hd__a221o_1 _2009_ (.A1(\dataMemory[24][6] ),
    .A2(net171),
    .B1(net140),
    .B2(\dataMemory[25][6] ),
    .C1(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__a211o_1 _2010_ (.A1(\dataMemory[26][6] ),
    .A2(net155),
    .B1(_1182_),
    .C1(net213),
    .X(_1183_));
 sky130_fd_sc_hd__mux4_1 _2011_ (.A0(\dataMemory[28][6] ),
    .A1(\dataMemory[29][6] ),
    .A2(\dataMemory[30][6] ),
    .A3(\dataMemory[31][6] ),
    .S0(net282),
    .S1(net244),
    .X(_1184_));
 sky130_fd_sc_hd__and3_1 _2012_ (.A(net282),
    .B(net244),
    .C(\dataMemory[7][6] ),
    .X(_1185_));
 sky130_fd_sc_hd__a221o_1 _2013_ (.A1(\dataMemory[6][6] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[5][6] ),
    .C1(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__a211o_1 _2014_ (.A1(\dataMemory[4][6] ),
    .A2(net171),
    .B1(_1186_),
    .C1(net189),
    .X(_1187_));
 sky130_fd_sc_hd__and3_1 _2015_ (.A(net282),
    .B(net244),
    .C(\dataMemory[3][6] ),
    .X(_1188_));
 sky130_fd_sc_hd__a221o_1 _2016_ (.A1(\dataMemory[2][6] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[1][6] ),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__a211o_1 _2017_ (.A1(\dataMemory[0][6] ),
    .A2(net171),
    .B1(_1189_),
    .C1(net213),
    .X(_1190_));
 sky130_fd_sc_hd__and3_1 _2018_ (.A(net282),
    .B(net244),
    .C(\dataMemory[11][6] ),
    .X(_1191_));
 sky130_fd_sc_hd__a221o_1 _2019_ (.A1(\dataMemory[8][6] ),
    .A2(net171),
    .B1(net140),
    .B2(\dataMemory[9][6] ),
    .C1(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__a211o_1 _2020_ (.A1(\dataMemory[10][6] ),
    .A2(net155),
    .B1(_1192_),
    .C1(net213),
    .X(_1193_));
 sky130_fd_sc_hd__mux4_1 _2021_ (.A0(\dataMemory[12][6] ),
    .A1(\dataMemory[13][6] ),
    .A2(\dataMemory[14][6] ),
    .A3(\dataMemory[15][6] ),
    .S0(net282),
    .S1(net244),
    .X(_1194_));
 sky130_fd_sc_hd__o21a_1 _2022_ (.A1(net189),
    .A2(_1194_),
    .B1(net207),
    .X(_1195_));
 sky130_fd_sc_hd__a32o_1 _2023_ (.A1(net184),
    .A2(_1187_),
    .A3(_1190_),
    .B1(_1193_),
    .B2(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__o21a_1 _2024_ (.A1(net189),
    .A2(_1184_),
    .B1(net207),
    .X(_1197_));
 sky130_fd_sc_hd__a32o_1 _2025_ (.A1(net184),
    .A2(_1177_),
    .A3(_1180_),
    .B1(_1183_),
    .B2(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_4 _2026_ (.A0(_1196_),
    .A1(_1198_),
    .S(net203),
    .X(net68));
 sky130_fd_sc_hd__and3_1 _2027_ (.A(net283),
    .B(net245),
    .C(\dataMemory[23][7] ),
    .X(_1199_));
 sky130_fd_sc_hd__a221o_1 _2028_ (.A1(\dataMemory[22][7] ),
    .A2(net155),
    .B1(net142),
    .B2(\dataMemory[21][7] ),
    .C1(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__a211o_1 _2029_ (.A1(\dataMemory[20][7] ),
    .A2(net173),
    .B1(_1200_),
    .C1(net189),
    .X(_1201_));
 sky130_fd_sc_hd__and3_1 _2030_ (.A(net283),
    .B(net245),
    .C(\dataMemory[19][7] ),
    .X(_1202_));
 sky130_fd_sc_hd__a221o_1 _2031_ (.A1(\dataMemory[18][7] ),
    .A2(net155),
    .B1(net142),
    .B2(\dataMemory[17][7] ),
    .C1(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__a211o_1 _2032_ (.A1(\dataMemory[16][7] ),
    .A2(net173),
    .B1(_1203_),
    .C1(net213),
    .X(_1204_));
 sky130_fd_sc_hd__and3_1 _2033_ (.A(net283),
    .B(net245),
    .C(\dataMemory[27][7] ),
    .X(_1205_));
 sky130_fd_sc_hd__a221o_1 _2034_ (.A1(\dataMemory[24][7] ),
    .A2(net173),
    .B1(net140),
    .B2(\dataMemory[25][7] ),
    .C1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__a211o_1 _2035_ (.A1(\dataMemory[26][7] ),
    .A2(net157),
    .B1(_1206_),
    .C1(net213),
    .X(_1207_));
 sky130_fd_sc_hd__mux4_1 _2036_ (.A0(\dataMemory[28][7] ),
    .A1(\dataMemory[29][7] ),
    .A2(\dataMemory[30][7] ),
    .A3(\dataMemory[31][7] ),
    .S0(net283),
    .S1(net245),
    .X(_1208_));
 sky130_fd_sc_hd__and3_1 _2037_ (.A(net283),
    .B(net245),
    .C(\dataMemory[7][7] ),
    .X(_1209_));
 sky130_fd_sc_hd__a221o_1 _2038_ (.A1(\dataMemory[6][7] ),
    .A2(net157),
    .B1(net140),
    .B2(\dataMemory[5][7] ),
    .C1(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__a211o_1 _2039_ (.A1(\dataMemory[4][7] ),
    .A2(net171),
    .B1(_1210_),
    .C1(net189),
    .X(_1211_));
 sky130_fd_sc_hd__and3_1 _2040_ (.A(net283),
    .B(net245),
    .C(\dataMemory[3][7] ),
    .X(_1212_));
 sky130_fd_sc_hd__a221o_1 _2041_ (.A1(\dataMemory[2][7] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[1][7] ),
    .C1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__a211o_1 _2042_ (.A1(\dataMemory[0][7] ),
    .A2(net171),
    .B1(_1213_),
    .C1(net213),
    .X(_1214_));
 sky130_fd_sc_hd__and3_1 _2043_ (.A(net283),
    .B(net245),
    .C(\dataMemory[11][7] ),
    .X(_1215_));
 sky130_fd_sc_hd__a221o_1 _2044_ (.A1(\dataMemory[8][7] ),
    .A2(net171),
    .B1(net140),
    .B2(\dataMemory[9][7] ),
    .C1(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__a211o_1 _2045_ (.A1(\dataMemory[10][7] ),
    .A2(net155),
    .B1(_1216_),
    .C1(net213),
    .X(_1217_));
 sky130_fd_sc_hd__mux4_1 _2046_ (.A0(\dataMemory[12][7] ),
    .A1(\dataMemory[13][7] ),
    .A2(\dataMemory[14][7] ),
    .A3(\dataMemory[15][7] ),
    .S0(net283),
    .S1(net245),
    .X(_1218_));
 sky130_fd_sc_hd__o21a_1 _2047_ (.A1(net189),
    .A2(_1218_),
    .B1(net207),
    .X(_1219_));
 sky130_fd_sc_hd__a32o_1 _2048_ (.A1(net184),
    .A2(_1211_),
    .A3(_1214_),
    .B1(_1217_),
    .B2(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__o21a_1 _2049_ (.A1(net189),
    .A2(_1208_),
    .B1(net207),
    .X(_1221_));
 sky130_fd_sc_hd__a32o_1 _2050_ (.A1(net184),
    .A2(_1201_),
    .A3(_1204_),
    .B1(_1207_),
    .B2(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__mux2_4 _2051_ (.A0(_1220_),
    .A1(_1222_),
    .S(net203),
    .X(net69));
 sky130_fd_sc_hd__and3_1 _2052_ (.A(net280),
    .B(net242),
    .C(\dataMemory[23][8] ),
    .X(_1223_));
 sky130_fd_sc_hd__a221o_1 _2053_ (.A1(\dataMemory[22][8] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[21][8] ),
    .C1(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__a211o_1 _2054_ (.A1(\dataMemory[20][8] ),
    .A2(net169),
    .B1(_1224_),
    .C1(net188),
    .X(_1225_));
 sky130_fd_sc_hd__and3_1 _2055_ (.A(net280),
    .B(net242),
    .C(\dataMemory[19][8] ),
    .X(_1226_));
 sky130_fd_sc_hd__a221o_1 _2056_ (.A1(\dataMemory[18][8] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[17][8] ),
    .C1(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__a211o_1 _2057_ (.A1(\dataMemory[16][8] ),
    .A2(net169),
    .B1(_1227_),
    .C1(net212),
    .X(_1228_));
 sky130_fd_sc_hd__and3_1 _2058_ (.A(net280),
    .B(net242),
    .C(\dataMemory[27][8] ),
    .X(_1229_));
 sky130_fd_sc_hd__a221o_1 _2059_ (.A1(\dataMemory[24][8] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[25][8] ),
    .C1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__a211o_1 _2060_ (.A1(\dataMemory[26][8] ),
    .A2(net153),
    .B1(_1230_),
    .C1(net212),
    .X(_1231_));
 sky130_fd_sc_hd__mux4_1 _2061_ (.A0(\dataMemory[28][8] ),
    .A1(\dataMemory[29][8] ),
    .A2(\dataMemory[30][8] ),
    .A3(\dataMemory[31][8] ),
    .S0(net280),
    .S1(net242),
    .X(_1232_));
 sky130_fd_sc_hd__and3_1 _2062_ (.A(net282),
    .B(net244),
    .C(\dataMemory[7][8] ),
    .X(_1233_));
 sky130_fd_sc_hd__a221o_1 _2063_ (.A1(\dataMemory[6][8] ),
    .A2(net152),
    .B1(net137),
    .B2(\dataMemory[5][8] ),
    .C1(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__a211o_1 _2064_ (.A1(\dataMemory[4][8] ),
    .A2(net171),
    .B1(_1234_),
    .C1(net196),
    .X(_1235_));
 sky130_fd_sc_hd__and3_1 _2065_ (.A(net283),
    .B(net245),
    .C(\dataMemory[3][8] ),
    .X(_1236_));
 sky130_fd_sc_hd__a221o_1 _2066_ (.A1(\dataMemory[2][8] ),
    .A2(net155),
    .B1(net140),
    .B2(\dataMemory[1][8] ),
    .C1(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__a211o_1 _2067_ (.A1(\dataMemory[0][8] ),
    .A2(net171),
    .B1(_1237_),
    .C1(net213),
    .X(_1238_));
 sky130_fd_sc_hd__and3_1 _2068_ (.A(net283),
    .B(net248),
    .C(\dataMemory[11][8] ),
    .X(_1239_));
 sky130_fd_sc_hd__a221o_1 _2069_ (.A1(\dataMemory[8][8] ),
    .A2(net168),
    .B1(net137),
    .B2(\dataMemory[9][8] ),
    .C1(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__a211o_1 _2070_ (.A1(\dataMemory[10][8] ),
    .A2(net152),
    .B1(_1240_),
    .C1(net215),
    .X(_1241_));
 sky130_fd_sc_hd__mux4_1 _2071_ (.A0(\dataMemory[12][8] ),
    .A1(\dataMemory[13][8] ),
    .A2(\dataMemory[14][8] ),
    .A3(\dataMemory[15][8] ),
    .S0(net284),
    .S1(net246),
    .X(_1242_));
 sky130_fd_sc_hd__o21a_1 _2072_ (.A1(net196),
    .A2(_1242_),
    .B1(net206),
    .X(_1243_));
 sky130_fd_sc_hd__a32o_1 _2073_ (.A1(net183),
    .A2(_1235_),
    .A3(_1238_),
    .B1(_1241_),
    .B2(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__o21a_1 _2074_ (.A1(net188),
    .A2(_1232_),
    .B1(net206),
    .X(_1245_));
 sky130_fd_sc_hd__a32o_1 _2075_ (.A1(net183),
    .A2(_1225_),
    .A3(_1228_),
    .B1(_1231_),
    .B2(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_4 _2076_ (.A0(_1244_),
    .A1(_1246_),
    .S(net203),
    .X(net70));
 sky130_fd_sc_hd__and3_1 _2077_ (.A(net280),
    .B(net242),
    .C(\dataMemory[23][9] ),
    .X(_1247_));
 sky130_fd_sc_hd__a221o_1 _2078_ (.A1(\dataMemory[22][9] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[21][9] ),
    .C1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__a211o_1 _2079_ (.A1(\dataMemory[20][9] ),
    .A2(net169),
    .B1(_1248_),
    .C1(net188),
    .X(_1249_));
 sky130_fd_sc_hd__and3_1 _2080_ (.A(net280),
    .B(net242),
    .C(\dataMemory[19][9] ),
    .X(_1250_));
 sky130_fd_sc_hd__a221o_1 _2081_ (.A1(\dataMemory[18][9] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[17][9] ),
    .C1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__a211o_1 _2082_ (.A1(\dataMemory[16][9] ),
    .A2(net169),
    .B1(_1251_),
    .C1(net212),
    .X(_1252_));
 sky130_fd_sc_hd__and3_1 _2083_ (.A(net280),
    .B(net242),
    .C(\dataMemory[27][9] ),
    .X(_1253_));
 sky130_fd_sc_hd__a221o_1 _2084_ (.A1(\dataMemory[24][9] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[25][9] ),
    .C1(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__a211o_1 _2085_ (.A1(\dataMemory[26][9] ),
    .A2(net153),
    .B1(_1254_),
    .C1(net212),
    .X(_1255_));
 sky130_fd_sc_hd__mux4_1 _2086_ (.A0(\dataMemory[28][9] ),
    .A1(\dataMemory[29][9] ),
    .A2(\dataMemory[30][9] ),
    .A3(\dataMemory[31][9] ),
    .S0(net280),
    .S1(net242),
    .X(_1256_));
 sky130_fd_sc_hd__and3_1 _2087_ (.A(net281),
    .B(net243),
    .C(\dataMemory[7][9] ),
    .X(_1257_));
 sky130_fd_sc_hd__a221o_1 _2088_ (.A1(\dataMemory[6][9] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[5][9] ),
    .C1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__a211o_1 _2089_ (.A1(\dataMemory[4][9] ),
    .A2(net170),
    .B1(_1258_),
    .C1(net188),
    .X(_1259_));
 sky130_fd_sc_hd__and3_1 _2090_ (.A(net281),
    .B(net243),
    .C(\dataMemory[3][9] ),
    .X(_1260_));
 sky130_fd_sc_hd__a221o_1 _2091_ (.A1(\dataMemory[2][9] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[1][9] ),
    .C1(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__a211o_1 _2092_ (.A1(\dataMemory[0][9] ),
    .A2(net170),
    .B1(_1261_),
    .C1(net212),
    .X(_1262_));
 sky130_fd_sc_hd__and3_1 _2093_ (.A(net281),
    .B(net243),
    .C(\dataMemory[11][9] ),
    .X(_1263_));
 sky130_fd_sc_hd__a221o_1 _2094_ (.A1(\dataMemory[8][9] ),
    .A2(net170),
    .B1(net138),
    .B2(\dataMemory[9][9] ),
    .C1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__a211o_1 _2095_ (.A1(\dataMemory[10][9] ),
    .A2(net154),
    .B1(_1264_),
    .C1(net212),
    .X(_1265_));
 sky130_fd_sc_hd__mux4_1 _2096_ (.A0(\dataMemory[12][9] ),
    .A1(\dataMemory[13][9] ),
    .A2(\dataMemory[14][9] ),
    .A3(\dataMemory[15][9] ),
    .S0(net281),
    .S1(net243),
    .X(_1266_));
 sky130_fd_sc_hd__o21a_1 _2097_ (.A1(net188),
    .A2(_1266_),
    .B1(net206),
    .X(_1267_));
 sky130_fd_sc_hd__a32o_1 _2098_ (.A1(net183),
    .A2(_1259_),
    .A3(_1262_),
    .B1(_1265_),
    .B2(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__o21a_1 _2099_ (.A1(net188),
    .A2(_1256_),
    .B1(net206),
    .X(_1269_));
 sky130_fd_sc_hd__a32o_1 _2100_ (.A1(net183),
    .A2(_1249_),
    .A3(_1252_),
    .B1(_1255_),
    .B2(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_4 _2101_ (.A0(_1268_),
    .A1(_1270_),
    .S(net203),
    .X(net71));
 sky130_fd_sc_hd__and3_1 _2102_ (.A(net285),
    .B(net247),
    .C(\dataMemory[23][10] ),
    .X(_1271_));
 sky130_fd_sc_hd__a221o_1 _2103_ (.A1(\dataMemory[22][10] ),
    .A2(net157),
    .B1(net142),
    .B2(\dataMemory[21][10] ),
    .C1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__a211o_1 _2104_ (.A1(\dataMemory[20][10] ),
    .A2(net173),
    .B1(_1272_),
    .C1(net190),
    .X(_1273_));
 sky130_fd_sc_hd__and3_1 _2105_ (.A(net285),
    .B(net247),
    .C(\dataMemory[19][10] ),
    .X(_1274_));
 sky130_fd_sc_hd__a221o_1 _2106_ (.A1(\dataMemory[18][10] ),
    .A2(net157),
    .B1(net142),
    .B2(\dataMemory[17][10] ),
    .C1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__a211o_1 _2107_ (.A1(\dataMemory[16][10] ),
    .A2(net173),
    .B1(_1275_),
    .C1(net213),
    .X(_1276_));
 sky130_fd_sc_hd__and3_1 _2108_ (.A(net283),
    .B(net245),
    .C(\dataMemory[27][10] ),
    .X(_1277_));
 sky130_fd_sc_hd__a221o_1 _2109_ (.A1(\dataMemory[24][10] ),
    .A2(net173),
    .B1(net142),
    .B2(\dataMemory[25][10] ),
    .C1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__a211o_1 _2110_ (.A1(\dataMemory[26][10] ),
    .A2(net157),
    .B1(_1278_),
    .C1(net213),
    .X(_1279_));
 sky130_fd_sc_hd__mux4_1 _2111_ (.A0(\dataMemory[28][10] ),
    .A1(\dataMemory[29][10] ),
    .A2(\dataMemory[30][10] ),
    .A3(\dataMemory[31][10] ),
    .S0(net285),
    .S1(net247),
    .X(_1280_));
 sky130_fd_sc_hd__and3_1 _2112_ (.A(net287),
    .B(net245),
    .C(\dataMemory[7][10] ),
    .X(_1281_));
 sky130_fd_sc_hd__a221o_1 _2113_ (.A1(\dataMemory[6][10] ),
    .A2(net157),
    .B1(net142),
    .B2(\dataMemory[5][10] ),
    .C1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__a211o_1 _2114_ (.A1(\dataMemory[4][10] ),
    .A2(net173),
    .B1(_1282_),
    .C1(net189),
    .X(_1283_));
 sky130_fd_sc_hd__and3_1 _2115_ (.A(net283),
    .B(net245),
    .C(\dataMemory[3][10] ),
    .X(_1284_));
 sky130_fd_sc_hd__a221o_1 _2116_ (.A1(\dataMemory[2][10] ),
    .A2(net157),
    .B1(net142),
    .B2(\dataMemory[1][10] ),
    .C1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__a211o_1 _2117_ (.A1(\dataMemory[0][10] ),
    .A2(net173),
    .B1(_1285_),
    .C1(net213),
    .X(_1286_));
 sky130_fd_sc_hd__and3_1 _2118_ (.A(net283),
    .B(net245),
    .C(\dataMemory[11][10] ),
    .X(_1287_));
 sky130_fd_sc_hd__a221o_1 _2119_ (.A1(\dataMemory[8][10] ),
    .A2(net173),
    .B1(net142),
    .B2(\dataMemory[9][10] ),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a211o_1 _2120_ (.A1(\dataMemory[10][10] ),
    .A2(net155),
    .B1(_1288_),
    .C1(net213),
    .X(_1289_));
 sky130_fd_sc_hd__mux4_1 _2121_ (.A0(\dataMemory[12][10] ),
    .A1(\dataMemory[13][10] ),
    .A2(\dataMemory[14][10] ),
    .A3(\dataMemory[15][10] ),
    .S0(net283),
    .S1(net245),
    .X(_1290_));
 sky130_fd_sc_hd__o21a_1 _2122_ (.A1(net189),
    .A2(_1290_),
    .B1(net207),
    .X(_1291_));
 sky130_fd_sc_hd__a32o_1 _2123_ (.A1(net184),
    .A2(_1283_),
    .A3(_1286_),
    .B1(_1289_),
    .B2(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__o21a_1 _2124_ (.A1(net189),
    .A2(_1280_),
    .B1(net207),
    .X(_1293_));
 sky130_fd_sc_hd__a32o_1 _2125_ (.A1(net184),
    .A2(_1273_),
    .A3(_1276_),
    .B1(_1279_),
    .B2(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_4 _2126_ (.A0(_1292_),
    .A1(_1294_),
    .S(net203),
    .X(net41));
 sky130_fd_sc_hd__and3_1 _2127_ (.A(net287),
    .B(net249),
    .C(\dataMemory[23][11] ),
    .X(_1295_));
 sky130_fd_sc_hd__a221o_1 _2128_ (.A1(\dataMemory[22][11] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[21][11] ),
    .C1(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__a211o_1 _2129_ (.A1(\dataMemory[20][11] ),
    .A2(net174),
    .B1(_1296_),
    .C1(net191),
    .X(_1297_));
 sky130_fd_sc_hd__and3_1 _2130_ (.A(net287),
    .B(net249),
    .C(\dataMemory[19][11] ),
    .X(_1298_));
 sky130_fd_sc_hd__a221o_1 _2131_ (.A1(\dataMemory[18][11] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[17][11] ),
    .C1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__a211o_1 _2132_ (.A1(\dataMemory[16][11] ),
    .A2(net175),
    .B1(_1299_),
    .C1(net216),
    .X(_1300_));
 sky130_fd_sc_hd__and3_1 _2133_ (.A(net287),
    .B(net249),
    .C(\dataMemory[27][11] ),
    .X(_1301_));
 sky130_fd_sc_hd__a221o_1 _2134_ (.A1(\dataMemory[24][11] ),
    .A2(net174),
    .B1(net143),
    .B2(\dataMemory[25][11] ),
    .C1(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__a211o_1 _2135_ (.A1(\dataMemory[26][11] ),
    .A2(net158),
    .B1(_1302_),
    .C1(net216),
    .X(_1303_));
 sky130_fd_sc_hd__mux4_1 _2136_ (.A0(\dataMemory[28][11] ),
    .A1(\dataMemory[29][11] ),
    .A2(\dataMemory[30][11] ),
    .A3(\dataMemory[31][11] ),
    .S0(net287),
    .S1(net249),
    .X(_1304_));
 sky130_fd_sc_hd__and3_1 _2137_ (.A(net291),
    .B(net253),
    .C(\dataMemory[7][11] ),
    .X(_1305_));
 sky130_fd_sc_hd__a221o_1 _2138_ (.A1(\dataMemory[6][11] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[5][11] ),
    .C1(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__a211o_1 _2139_ (.A1(\dataMemory[4][11] ),
    .A2(net179),
    .B1(_1306_),
    .C1(net193),
    .X(_1307_));
 sky130_fd_sc_hd__and3_1 _2140_ (.A(net288),
    .B(net249),
    .C(\dataMemory[3][11] ),
    .X(_1308_));
 sky130_fd_sc_hd__a221o_1 _2141_ (.A1(\dataMemory[2][11] ),
    .A2(net159),
    .B1(net145),
    .B2(\dataMemory[1][11] ),
    .C1(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__a211o_1 _2142_ (.A1(\dataMemory[0][11] ),
    .A2(net179),
    .B1(_1309_),
    .C1(net218),
    .X(_1310_));
 sky130_fd_sc_hd__and3_1 _2143_ (.A(net288),
    .B(net250),
    .C(\dataMemory[11][11] ),
    .X(_1311_));
 sky130_fd_sc_hd__a221o_1 _2144_ (.A1(\dataMemory[8][11] ),
    .A2(net175),
    .B1(net145),
    .B2(\dataMemory[9][11] ),
    .C1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__a211o_1 _2145_ (.A1(\dataMemory[10][11] ),
    .A2(net159),
    .B1(_1312_),
    .C1(net218),
    .X(_1313_));
 sky130_fd_sc_hd__mux4_1 _2146_ (.A0(\dataMemory[12][11] ),
    .A1(\dataMemory[13][11] ),
    .A2(\dataMemory[14][11] ),
    .A3(\dataMemory[15][11] ),
    .S0(net288),
    .S1(net250),
    .X(_1314_));
 sky130_fd_sc_hd__o21a_1 _2147_ (.A1(net191),
    .A2(_1314_),
    .B1(net208),
    .X(_1315_));
 sky130_fd_sc_hd__a32o_1 _2148_ (.A1(net185),
    .A2(_1307_),
    .A3(_1310_),
    .B1(_1313_),
    .B2(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__o21a_1 _2149_ (.A1(net191),
    .A2(_1304_),
    .B1(net209),
    .X(_1317_));
 sky130_fd_sc_hd__a32o_1 _2150_ (.A1(net186),
    .A2(_1297_),
    .A3(_1300_),
    .B1(_1303_),
    .B2(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_2 _2151_ (.A0(_1316_),
    .A1(_1318_),
    .S(net204),
    .X(net42));
 sky130_fd_sc_hd__and3_1 _2152_ (.A(net287),
    .B(net249),
    .C(\dataMemory[23][12] ),
    .X(_1319_));
 sky130_fd_sc_hd__a221o_1 _2153_ (.A1(\dataMemory[22][12] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[21][12] ),
    .C1(_1319_),
    .X(_1320_));
 sky130_fd_sc_hd__a211o_1 _2154_ (.A1(\dataMemory[20][12] ),
    .A2(net174),
    .B1(_1320_),
    .C1(net191),
    .X(_1321_));
 sky130_fd_sc_hd__and3_1 _2155_ (.A(net287),
    .B(net249),
    .C(\dataMemory[19][12] ),
    .X(_1322_));
 sky130_fd_sc_hd__a221o_1 _2156_ (.A1(\dataMemory[18][12] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[17][12] ),
    .C1(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__a211o_1 _2157_ (.A1(\dataMemory[16][12] ),
    .A2(net174),
    .B1(_1323_),
    .C1(net216),
    .X(_1324_));
 sky130_fd_sc_hd__and3_1 _2158_ (.A(net283),
    .B(net245),
    .C(\dataMemory[27][12] ),
    .X(_1325_));
 sky130_fd_sc_hd__a221o_1 _2159_ (.A1(\dataMemory[24][12] ),
    .A2(net171),
    .B1(net140),
    .B2(\dataMemory[25][12] ),
    .C1(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__a211o_1 _2160_ (.A1(\dataMemory[26][12] ),
    .A2(net155),
    .B1(_1326_),
    .C1(net213),
    .X(_1327_));
 sky130_fd_sc_hd__mux4_1 _2161_ (.A0(\dataMemory[28][12] ),
    .A1(\dataMemory[29][12] ),
    .A2(\dataMemory[30][12] ),
    .A3(\dataMemory[31][12] ),
    .S0(net287),
    .S1(net249),
    .X(_1328_));
 sky130_fd_sc_hd__and3_1 _2162_ (.A(net287),
    .B(net249),
    .C(\dataMemory[7][12] ),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _2163_ (.A1(\dataMemory[6][12] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[5][12] ),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__a211o_1 _2164_ (.A1(\dataMemory[4][12] ),
    .A2(net174),
    .B1(_1330_),
    .C1(net191),
    .X(_1331_));
 sky130_fd_sc_hd__and3_1 _2165_ (.A(net287),
    .B(net249),
    .C(\dataMemory[3][12] ),
    .X(_1332_));
 sky130_fd_sc_hd__a221o_1 _2166_ (.A1(\dataMemory[2][12] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[1][12] ),
    .C1(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__a211o_1 _2167_ (.A1(\dataMemory[0][12] ),
    .A2(net174),
    .B1(_1333_),
    .C1(net216),
    .X(_1334_));
 sky130_fd_sc_hd__and3_1 _2168_ (.A(net287),
    .B(net248),
    .C(\dataMemory[11][12] ),
    .X(_1335_));
 sky130_fd_sc_hd__a221o_1 _2169_ (.A1(\dataMemory[8][12] ),
    .A2(net174),
    .B1(net140),
    .B2(\dataMemory[9][12] ),
    .C1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__a211o_1 _2170_ (.A1(\dataMemory[10][12] ),
    .A2(net158),
    .B1(_1336_),
    .C1(net216),
    .X(_1337_));
 sky130_fd_sc_hd__mux4_1 _2171_ (.A0(\dataMemory[12][12] ),
    .A1(\dataMemory[13][12] ),
    .A2(\dataMemory[14][12] ),
    .A3(\dataMemory[15][12] ),
    .S0(net287),
    .S1(net249),
    .X(_1338_));
 sky130_fd_sc_hd__o21a_1 _2172_ (.A1(net191),
    .A2(_1338_),
    .B1(net209),
    .X(_1339_));
 sky130_fd_sc_hd__a32o_1 _2173_ (.A1(net186),
    .A2(_1331_),
    .A3(_1334_),
    .B1(_1337_),
    .B2(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__o21a_1 _2174_ (.A1(net191),
    .A2(_1328_),
    .B1(net209),
    .X(_1341_));
 sky130_fd_sc_hd__a32o_1 _2175_ (.A1(net186),
    .A2(_1321_),
    .A3(_1324_),
    .B1(_1327_),
    .B2(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__mux2_4 _2176_ (.A0(_1340_),
    .A1(_1342_),
    .S(net203),
    .X(net43));
 sky130_fd_sc_hd__and3_1 _2177_ (.A(net281),
    .B(net243),
    .C(\dataMemory[23][13] ),
    .X(_1343_));
 sky130_fd_sc_hd__a221o_1 _2178_ (.A1(\dataMemory[22][13] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[21][13] ),
    .C1(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__a211o_1 _2179_ (.A1(\dataMemory[20][13] ),
    .A2(net170),
    .B1(_1344_),
    .C1(net188),
    .X(_1345_));
 sky130_fd_sc_hd__and3_1 _2180_ (.A(net281),
    .B(net243),
    .C(\dataMemory[19][13] ),
    .X(_1346_));
 sky130_fd_sc_hd__a221o_1 _2181_ (.A1(\dataMemory[18][13] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[17][13] ),
    .C1(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a211o_1 _2182_ (.A1(\dataMemory[16][13] ),
    .A2(net170),
    .B1(_1347_),
    .C1(net212),
    .X(_1348_));
 sky130_fd_sc_hd__and3_1 _2183_ (.A(net280),
    .B(net242),
    .C(\dataMemory[27][13] ),
    .X(_1349_));
 sky130_fd_sc_hd__a221o_1 _2184_ (.A1(\dataMemory[24][13] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[25][13] ),
    .C1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__a211o_1 _2185_ (.A1(\dataMemory[26][13] ),
    .A2(net153),
    .B1(_1350_),
    .C1(net212),
    .X(_1351_));
 sky130_fd_sc_hd__mux4_1 _2186_ (.A0(\dataMemory[28][13] ),
    .A1(\dataMemory[29][13] ),
    .A2(\dataMemory[30][13] ),
    .A3(\dataMemory[31][13] ),
    .S0(net281),
    .S1(net243),
    .X(_1352_));
 sky130_fd_sc_hd__and3_1 _2187_ (.A(net284),
    .B(net246),
    .C(\dataMemory[7][13] ),
    .X(_1353_));
 sky130_fd_sc_hd__a221o_1 _2188_ (.A1(\dataMemory[6][13] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[5][13] ),
    .C1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__a211o_1 _2189_ (.A1(\dataMemory[4][13] ),
    .A2(net172),
    .B1(_1354_),
    .C1(net190),
    .X(_1355_));
 sky130_fd_sc_hd__and3_1 _2190_ (.A(net284),
    .B(net246),
    .C(\dataMemory[3][13] ),
    .X(_1356_));
 sky130_fd_sc_hd__a221o_1 _2191_ (.A1(\dataMemory[2][13] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[1][13] ),
    .C1(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__a211o_1 _2192_ (.A1(\dataMemory[0][13] ),
    .A2(net172),
    .B1(_1357_),
    .C1(net214),
    .X(_1358_));
 sky130_fd_sc_hd__and3_1 _2193_ (.A(net284),
    .B(net246),
    .C(\dataMemory[11][13] ),
    .X(_1359_));
 sky130_fd_sc_hd__a221o_1 _2194_ (.A1(\dataMemory[8][13] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[9][13] ),
    .C1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__a211o_1 _2195_ (.A1(\dataMemory[10][13] ),
    .A2(net156),
    .B1(_1360_),
    .C1(net214),
    .X(_1361_));
 sky130_fd_sc_hd__mux4_1 _2196_ (.A0(\dataMemory[12][13] ),
    .A1(\dataMemory[13][13] ),
    .A2(\dataMemory[14][13] ),
    .A3(\dataMemory[15][13] ),
    .S0(net284),
    .S1(net246),
    .X(_1362_));
 sky130_fd_sc_hd__o21a_1 _2197_ (.A1(net190),
    .A2(_1362_),
    .B1(net207),
    .X(_1363_));
 sky130_fd_sc_hd__a32o_1 _2198_ (.A1(_1025_),
    .A2(_1355_),
    .A3(_1358_),
    .B1(_1361_),
    .B2(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__o21a_1 _2199_ (.A1(net188),
    .A2(_1352_),
    .B1(net206),
    .X(_1365_));
 sky130_fd_sc_hd__a32o_1 _2200_ (.A1(net183),
    .A2(_1345_),
    .A3(_1348_),
    .B1(_1351_),
    .B2(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_4 _2201_ (.A0(_1364_),
    .A1(_1366_),
    .S(net203),
    .X(net44));
 sky130_fd_sc_hd__and3_1 _2202_ (.A(net284),
    .B(net246),
    .C(\dataMemory[23][14] ),
    .X(_1367_));
 sky130_fd_sc_hd__a221o_1 _2203_ (.A1(\dataMemory[22][14] ),
    .A2(net154),
    .B1(net139),
    .B2(\dataMemory[21][14] ),
    .C1(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__a211o_1 _2204_ (.A1(\dataMemory[20][14] ),
    .A2(net170),
    .B1(_1368_),
    .C1(net188),
    .X(_1369_));
 sky130_fd_sc_hd__and3_1 _2205_ (.A(net284),
    .B(net246),
    .C(\dataMemory[19][14] ),
    .X(_1370_));
 sky130_fd_sc_hd__a221o_1 _2206_ (.A1(\dataMemory[18][14] ),
    .A2(net153),
    .B1(net139),
    .B2(\dataMemory[17][14] ),
    .C1(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__a211o_1 _2207_ (.A1(\dataMemory[16][14] ),
    .A2(net169),
    .B1(_1371_),
    .C1(net212),
    .X(_1372_));
 sky130_fd_sc_hd__and3_1 _2208_ (.A(net281),
    .B(net243),
    .C(\dataMemory[27][14] ),
    .X(_1373_));
 sky130_fd_sc_hd__a221o_1 _2209_ (.A1(\dataMemory[24][14] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[25][14] ),
    .C1(_1373_),
    .X(_1374_));
 sky130_fd_sc_hd__a211o_1 _2210_ (.A1(\dataMemory[26][14] ),
    .A2(net153),
    .B1(_1374_),
    .C1(net212),
    .X(_1375_));
 sky130_fd_sc_hd__mux4_1 _2211_ (.A0(\dataMemory[28][14] ),
    .A1(\dataMemory[29][14] ),
    .A2(\dataMemory[30][14] ),
    .A3(\dataMemory[31][14] ),
    .S0(net281),
    .S1(net243),
    .X(_1376_));
 sky130_fd_sc_hd__and3_1 _2212_ (.A(net284),
    .B(net246),
    .C(\dataMemory[7][14] ),
    .X(_1377_));
 sky130_fd_sc_hd__a221o_1 _2213_ (.A1(\dataMemory[6][14] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[5][14] ),
    .C1(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__a211o_1 _2214_ (.A1(\dataMemory[4][14] ),
    .A2(net169),
    .B1(_1378_),
    .C1(net188),
    .X(_1379_));
 sky130_fd_sc_hd__and3_1 _2215_ (.A(net284),
    .B(net246),
    .C(\dataMemory[3][14] ),
    .X(_1380_));
 sky130_fd_sc_hd__a221o_1 _2216_ (.A1(\dataMemory[2][14] ),
    .A2(net153),
    .B1(net138),
    .B2(\dataMemory[1][14] ),
    .C1(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__a211o_1 _2217_ (.A1(\dataMemory[0][14] ),
    .A2(net169),
    .B1(_1381_),
    .C1(net212),
    .X(_1382_));
 sky130_fd_sc_hd__and3_1 _2218_ (.A(net281),
    .B(net243),
    .C(\dataMemory[11][14] ),
    .X(_1383_));
 sky130_fd_sc_hd__a221o_1 _2219_ (.A1(\dataMemory[8][14] ),
    .A2(net169),
    .B1(net138),
    .B2(\dataMemory[9][14] ),
    .C1(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__a211o_1 _2220_ (.A1(\dataMemory[10][14] ),
    .A2(net153),
    .B1(_1384_),
    .C1(net215),
    .X(_1385_));
 sky130_fd_sc_hd__mux4_1 _2221_ (.A0(\dataMemory[12][14] ),
    .A1(\dataMemory[13][14] ),
    .A2(\dataMemory[14][14] ),
    .A3(\dataMemory[15][14] ),
    .S0(net281),
    .S1(net243),
    .X(_1386_));
 sky130_fd_sc_hd__o21a_1 _2222_ (.A1(net188),
    .A2(_1386_),
    .B1(net207),
    .X(_1387_));
 sky130_fd_sc_hd__a32o_1 _2223_ (.A1(net183),
    .A2(_1379_),
    .A3(_1382_),
    .B1(_1385_),
    .B2(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__o21a_1 _2224_ (.A1(net188),
    .A2(_1376_),
    .B1(net207),
    .X(_1389_));
 sky130_fd_sc_hd__a32o_1 _2225_ (.A1(net183),
    .A2(_1369_),
    .A3(_1372_),
    .B1(_1375_),
    .B2(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_4 _2226_ (.A0(_1388_),
    .A1(_1390_),
    .S(net203),
    .X(net45));
 sky130_fd_sc_hd__and3_1 _2227_ (.A(net287),
    .B(net249),
    .C(\dataMemory[23][15] ),
    .X(_1391_));
 sky130_fd_sc_hd__a221o_1 _2228_ (.A1(\dataMemory[22][15] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[21][15] ),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__a211o_1 _2229_ (.A1(\dataMemory[20][15] ),
    .A2(net174),
    .B1(_1392_),
    .C1(net191),
    .X(_1393_));
 sky130_fd_sc_hd__and3_1 _2230_ (.A(net289),
    .B(net252),
    .C(\dataMemory[19][15] ),
    .X(_1394_));
 sky130_fd_sc_hd__a221o_1 _2231_ (.A1(\dataMemory[18][15] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[17][15] ),
    .C1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__a211o_1 _2232_ (.A1(\dataMemory[16][15] ),
    .A2(net176),
    .B1(_1395_),
    .C1(net216),
    .X(_1396_));
 sky130_fd_sc_hd__and3_1 _2233_ (.A(net287),
    .B(net249),
    .C(\dataMemory[27][15] ),
    .X(_1397_));
 sky130_fd_sc_hd__a221o_1 _2234_ (.A1(\dataMemory[24][15] ),
    .A2(net174),
    .B1(net143),
    .B2(\dataMemory[25][15] ),
    .C1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__a211o_1 _2235_ (.A1(\dataMemory[26][15] ),
    .A2(net158),
    .B1(_1398_),
    .C1(net216),
    .X(_1399_));
 sky130_fd_sc_hd__mux4_1 _2236_ (.A0(\dataMemory[28][15] ),
    .A1(\dataMemory[29][15] ),
    .A2(\dataMemory[30][15] ),
    .A3(\dataMemory[31][15] ),
    .S0(net289),
    .S1(net252),
    .X(_1400_));
 sky130_fd_sc_hd__and3_1 _2237_ (.A(net287),
    .B(net249),
    .C(\dataMemory[7][15] ),
    .X(_1401_));
 sky130_fd_sc_hd__a221o_1 _2238_ (.A1(\dataMemory[6][15] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[5][15] ),
    .C1(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__a211o_1 _2239_ (.A1(\dataMemory[4][15] ),
    .A2(net174),
    .B1(_1402_),
    .C1(net191),
    .X(_1403_));
 sky130_fd_sc_hd__and3_1 _2240_ (.A(net288),
    .B(net250),
    .C(\dataMemory[3][15] ),
    .X(_1404_));
 sky130_fd_sc_hd__a221o_1 _2241_ (.A1(\dataMemory[2][15] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[1][15] ),
    .C1(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__a211o_1 _2242_ (.A1(\dataMemory[0][15] ),
    .A2(net174),
    .B1(_1405_),
    .C1(net216),
    .X(_1406_));
 sky130_fd_sc_hd__and3_1 _2243_ (.A(net287),
    .B(net249),
    .C(\dataMemory[11][15] ),
    .X(_1407_));
 sky130_fd_sc_hd__a221o_1 _2244_ (.A1(\dataMemory[8][15] ),
    .A2(net174),
    .B1(net143),
    .B2(\dataMemory[9][15] ),
    .C1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__a211o_1 _2245_ (.A1(\dataMemory[10][15] ),
    .A2(net158),
    .B1(_1408_),
    .C1(net216),
    .X(_1409_));
 sky130_fd_sc_hd__mux4_1 _2246_ (.A0(\dataMemory[12][15] ),
    .A1(\dataMemory[13][15] ),
    .A2(\dataMemory[14][15] ),
    .A3(\dataMemory[15][15] ),
    .S0(net288),
    .S1(net249),
    .X(_1410_));
 sky130_fd_sc_hd__o21a_1 _2247_ (.A1(net191),
    .A2(_1410_),
    .B1(net209),
    .X(_1411_));
 sky130_fd_sc_hd__a32o_1 _2248_ (.A1(net186),
    .A2(_1403_),
    .A3(_1406_),
    .B1(_1409_),
    .B2(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__o21a_1 _2249_ (.A1(net192),
    .A2(_1400_),
    .B1(net209),
    .X(_1413_));
 sky130_fd_sc_hd__a32o_1 _2250_ (.A1(net186),
    .A2(_1393_),
    .A3(_1396_),
    .B1(_1399_),
    .B2(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_2 _2251_ (.A0(_1412_),
    .A1(_1414_),
    .S(net204),
    .X(net46));
 sky130_fd_sc_hd__and3_1 _2252_ (.A(net288),
    .B(net250),
    .C(\dataMemory[23][16] ),
    .X(_1415_));
 sky130_fd_sc_hd__a221o_1 _2253_ (.A1(\dataMemory[22][16] ),
    .A2(net159),
    .B1(net145),
    .B2(\dataMemory[21][16] ),
    .C1(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__a211o_1 _2254_ (.A1(\dataMemory[20][16] ),
    .A2(net175),
    .B1(_1416_),
    .C1(net191),
    .X(_1417_));
 sky130_fd_sc_hd__and3_1 _2255_ (.A(net288),
    .B(net250),
    .C(\dataMemory[19][16] ),
    .X(_1418_));
 sky130_fd_sc_hd__a221o_1 _2256_ (.A1(\dataMemory[18][16] ),
    .A2(net159),
    .B1(net145),
    .B2(\dataMemory[17][16] ),
    .C1(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__a211o_1 _2257_ (.A1(\dataMemory[16][16] ),
    .A2(net175),
    .B1(_1419_),
    .C1(net216),
    .X(_1420_));
 sky130_fd_sc_hd__and3_1 _2258_ (.A(net288),
    .B(net250),
    .C(\dataMemory[27][16] ),
    .X(_1421_));
 sky130_fd_sc_hd__a221o_1 _2259_ (.A1(\dataMemory[24][16] ),
    .A2(net175),
    .B1(net145),
    .B2(\dataMemory[25][16] ),
    .C1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__a211o_1 _2260_ (.A1(\dataMemory[26][16] ),
    .A2(net159),
    .B1(_1422_),
    .C1(net216),
    .X(_1423_));
 sky130_fd_sc_hd__mux4_1 _2261_ (.A0(\dataMemory[28][16] ),
    .A1(\dataMemory[29][16] ),
    .A2(\dataMemory[30][16] ),
    .A3(\dataMemory[31][16] ),
    .S0(net288),
    .S1(net250),
    .X(_1424_));
 sky130_fd_sc_hd__and3_1 _2262_ (.A(net292),
    .B(net254),
    .C(\dataMemory[7][16] ),
    .X(_1425_));
 sky130_fd_sc_hd__a221o_1 _2263_ (.A1(\dataMemory[6][16] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[5][16] ),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a211o_1 _2264_ (.A1(\dataMemory[4][16] ),
    .A2(net178),
    .B1(_1426_),
    .C1(net195),
    .X(_1427_));
 sky130_fd_sc_hd__and3_1 _2265_ (.A(net292),
    .B(net254),
    .C(\dataMemory[3][16] ),
    .X(_1428_));
 sky130_fd_sc_hd__a221o_1 _2266_ (.A1(\dataMemory[2][16] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[1][16] ),
    .C1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__a211o_1 _2267_ (.A1(\dataMemory[0][16] ),
    .A2(net178),
    .B1(_1429_),
    .C1(net218),
    .X(_1430_));
 sky130_fd_sc_hd__and3_1 _2268_ (.A(net292),
    .B(net254),
    .C(\dataMemory[11][16] ),
    .X(_1431_));
 sky130_fd_sc_hd__a221o_1 _2269_ (.A1(\dataMemory[8][16] ),
    .A2(net178),
    .B1(net147),
    .B2(\dataMemory[9][16] ),
    .C1(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__a211o_1 _2270_ (.A1(\dataMemory[10][16] ),
    .A2(net163),
    .B1(_1432_),
    .C1(net219),
    .X(_1433_));
 sky130_fd_sc_hd__mux4_1 _2271_ (.A0(\dataMemory[12][16] ),
    .A1(\dataMemory[13][16] ),
    .A2(\dataMemory[14][16] ),
    .A3(\dataMemory[15][16] ),
    .S0(net292),
    .S1(net254),
    .X(_1434_));
 sky130_fd_sc_hd__o21a_1 _2272_ (.A1(net195),
    .A2(_1434_),
    .B1(net208),
    .X(_1435_));
 sky130_fd_sc_hd__a32o_1 _2273_ (.A1(net185),
    .A2(_1427_),
    .A3(_1430_),
    .B1(_1433_),
    .B2(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__o21a_1 _2274_ (.A1(net191),
    .A2(_1424_),
    .B1(net209),
    .X(_1437_));
 sky130_fd_sc_hd__a32o_1 _2275_ (.A1(net186),
    .A2(_1417_),
    .A3(_1420_),
    .B1(_1423_),
    .B2(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__mux2_2 _2276_ (.A0(_1436_),
    .A1(_1438_),
    .S(net204),
    .X(net47));
 sky130_fd_sc_hd__and3_1 _2277_ (.A(net288),
    .B(net250),
    .C(\dataMemory[23][17] ),
    .X(_1439_));
 sky130_fd_sc_hd__a221o_1 _2278_ (.A1(\dataMemory[22][17] ),
    .A2(net159),
    .B1(net145),
    .B2(\dataMemory[21][17] ),
    .C1(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__a211o_1 _2279_ (.A1(\dataMemory[20][17] ),
    .A2(net174),
    .B1(_1440_),
    .C1(net191),
    .X(_1441_));
 sky130_fd_sc_hd__and3_1 _2280_ (.A(net288),
    .B(net250),
    .C(\dataMemory[19][17] ),
    .X(_1442_));
 sky130_fd_sc_hd__a221o_1 _2281_ (.A1(\dataMemory[18][17] ),
    .A2(net159),
    .B1(net143),
    .B2(\dataMemory[17][17] ),
    .C1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__a211o_1 _2282_ (.A1(\dataMemory[16][17] ),
    .A2(net174),
    .B1(_1443_),
    .C1(net216),
    .X(_1444_));
 sky130_fd_sc_hd__and3_1 _2283_ (.A(net288),
    .B(net250),
    .C(\dataMemory[27][17] ),
    .X(_1445_));
 sky130_fd_sc_hd__a221o_1 _2284_ (.A1(\dataMemory[24][17] ),
    .A2(net175),
    .B1(net145),
    .B2(\dataMemory[25][17] ),
    .C1(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__a211o_1 _2285_ (.A1(\dataMemory[26][17] ),
    .A2(net158),
    .B1(_1446_),
    .C1(net216),
    .X(_1447_));
 sky130_fd_sc_hd__mux4_1 _2286_ (.A0(\dataMemory[28][17] ),
    .A1(\dataMemory[29][17] ),
    .A2(\dataMemory[30][17] ),
    .A3(\dataMemory[31][17] ),
    .S0(net288),
    .S1(net250),
    .X(_1448_));
 sky130_fd_sc_hd__and3_1 _2287_ (.A(net292),
    .B(net254),
    .C(\dataMemory[7][17] ),
    .X(_1449_));
 sky130_fd_sc_hd__a221o_1 _2288_ (.A1(\dataMemory[6][17] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[5][17] ),
    .C1(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__a211o_1 _2289_ (.A1(\dataMemory[4][17] ),
    .A2(net178),
    .B1(_1450_),
    .C1(net195),
    .X(_1451_));
 sky130_fd_sc_hd__and3_1 _2290_ (.A(net292),
    .B(net254),
    .C(\dataMemory[3][17] ),
    .X(_1452_));
 sky130_fd_sc_hd__a221o_1 _2291_ (.A1(\dataMemory[2][17] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[1][17] ),
    .C1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__a211o_1 _2292_ (.A1(\dataMemory[0][17] ),
    .A2(net178),
    .B1(_1453_),
    .C1(net219),
    .X(_1454_));
 sky130_fd_sc_hd__and3_1 _2293_ (.A(net291),
    .B(net253),
    .C(\dataMemory[11][17] ),
    .X(_1455_));
 sky130_fd_sc_hd__a221o_1 _2294_ (.A1(\dataMemory[8][17] ),
    .A2(net178),
    .B1(net146),
    .B2(\dataMemory[9][17] ),
    .C1(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__a211o_1 _2295_ (.A1(\dataMemory[10][17] ),
    .A2(net163),
    .B1(_1456_),
    .C1(net219),
    .X(_1457_));
 sky130_fd_sc_hd__mux4_1 _2296_ (.A0(\dataMemory[12][17] ),
    .A1(\dataMemory[13][17] ),
    .A2(\dataMemory[14][17] ),
    .A3(\dataMemory[15][17] ),
    .S0(net291),
    .S1(net253),
    .X(_1458_));
 sky130_fd_sc_hd__o21a_1 _2297_ (.A1(net193),
    .A2(_1458_),
    .B1(net208),
    .X(_1459_));
 sky130_fd_sc_hd__a32o_1 _2298_ (.A1(net185),
    .A2(_1451_),
    .A3(_1454_),
    .B1(_1457_),
    .B2(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__o21a_1 _2299_ (.A1(net191),
    .A2(_1448_),
    .B1(net209),
    .X(_1461_));
 sky130_fd_sc_hd__a32o_1 _2300_ (.A1(net186),
    .A2(_1441_),
    .A3(_1444_),
    .B1(_1447_),
    .B2(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_2 _2301_ (.A0(_1460_),
    .A1(_1462_),
    .S(net204),
    .X(net48));
 sky130_fd_sc_hd__and3_1 _2302_ (.A(net289),
    .B(net252),
    .C(\dataMemory[23][18] ),
    .X(_1463_));
 sky130_fd_sc_hd__a221o_1 _2303_ (.A1(\dataMemory[22][18] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[21][18] ),
    .C1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__a211o_1 _2304_ (.A1(\dataMemory[20][18] ),
    .A2(net176),
    .B1(_1464_),
    .C1(net192),
    .X(_1465_));
 sky130_fd_sc_hd__and3_1 _2305_ (.A(net289),
    .B(net252),
    .C(\dataMemory[19][18] ),
    .X(_1466_));
 sky130_fd_sc_hd__a221o_1 _2306_ (.A1(\dataMemory[18][18] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[17][18] ),
    .C1(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__a211o_1 _2307_ (.A1(\dataMemory[16][18] ),
    .A2(net176),
    .B1(_1467_),
    .C1(net217),
    .X(_1468_));
 sky130_fd_sc_hd__and3_1 _2308_ (.A(net289),
    .B(net252),
    .C(\dataMemory[27][18] ),
    .X(_1469_));
 sky130_fd_sc_hd__a221o_1 _2309_ (.A1(\dataMemory[24][18] ),
    .A2(net176),
    .B1(net144),
    .B2(\dataMemory[25][18] ),
    .C1(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__a211o_1 _2310_ (.A1(\dataMemory[26][18] ),
    .A2(net160),
    .B1(_1470_),
    .C1(net217),
    .X(_1471_));
 sky130_fd_sc_hd__mux4_1 _2311_ (.A0(\dataMemory[28][18] ),
    .A1(\dataMemory[29][18] ),
    .A2(\dataMemory[30][18] ),
    .A3(\dataMemory[31][18] ),
    .S0(net289),
    .S1(net252),
    .X(_1472_));
 sky130_fd_sc_hd__and3_1 _2312_ (.A(net289),
    .B(net252),
    .C(\dataMemory[7][18] ),
    .X(_1473_));
 sky130_fd_sc_hd__a221o_1 _2313_ (.A1(\dataMemory[6][18] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[5][18] ),
    .C1(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__a211o_1 _2314_ (.A1(\dataMemory[4][18] ),
    .A2(net176),
    .B1(_1474_),
    .C1(net192),
    .X(_1475_));
 sky130_fd_sc_hd__and3_1 _2315_ (.A(net289),
    .B(net252),
    .C(\dataMemory[3][18] ),
    .X(_1476_));
 sky130_fd_sc_hd__a221o_1 _2316_ (.A1(\dataMemory[2][18] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[1][18] ),
    .C1(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__a211o_1 _2317_ (.A1(\dataMemory[0][18] ),
    .A2(net176),
    .B1(_1477_),
    .C1(net217),
    .X(_1478_));
 sky130_fd_sc_hd__and3_1 _2318_ (.A(net289),
    .B(net252),
    .C(\dataMemory[11][18] ),
    .X(_1479_));
 sky130_fd_sc_hd__a221o_1 _2319_ (.A1(\dataMemory[8][18] ),
    .A2(net176),
    .B1(net144),
    .B2(\dataMemory[9][18] ),
    .C1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__a211o_1 _2320_ (.A1(\dataMemory[10][18] ),
    .A2(net160),
    .B1(_1480_),
    .C1(net217),
    .X(_1481_));
 sky130_fd_sc_hd__mux4_1 _2321_ (.A0(\dataMemory[12][18] ),
    .A1(\dataMemory[13][18] ),
    .A2(\dataMemory[14][18] ),
    .A3(\dataMemory[15][18] ),
    .S0(net289),
    .S1(net252),
    .X(_1482_));
 sky130_fd_sc_hd__o21a_1 _2322_ (.A1(net192),
    .A2(_1482_),
    .B1(net209),
    .X(_1483_));
 sky130_fd_sc_hd__a32o_1 _2323_ (.A1(net186),
    .A2(_1475_),
    .A3(_1478_),
    .B1(_1481_),
    .B2(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__o21a_1 _2324_ (.A1(net192),
    .A2(_1472_),
    .B1(net209),
    .X(_1485_));
 sky130_fd_sc_hd__a32o_1 _2325_ (.A1(net186),
    .A2(_1465_),
    .A3(_1468_),
    .B1(_1471_),
    .B2(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_2 _2326_ (.A0(_1484_),
    .A1(_1486_),
    .S(net204),
    .X(net49));
 sky130_fd_sc_hd__and3_1 _2327_ (.A(net284),
    .B(net246),
    .C(\dataMemory[23][19] ),
    .X(_1487_));
 sky130_fd_sc_hd__a221o_1 _2328_ (.A1(\dataMemory[22][19] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[21][19] ),
    .C1(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__a211o_1 _2329_ (.A1(\dataMemory[20][19] ),
    .A2(net172),
    .B1(_1488_),
    .C1(net190),
    .X(_1489_));
 sky130_fd_sc_hd__and3_1 _2330_ (.A(net284),
    .B(net246),
    .C(\dataMemory[19][19] ),
    .X(_1490_));
 sky130_fd_sc_hd__a221o_1 _2331_ (.A1(\dataMemory[18][19] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[17][19] ),
    .C1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a211o_1 _2332_ (.A1(\dataMemory[16][19] ),
    .A2(net172),
    .B1(_1491_),
    .C1(net214),
    .X(_1492_));
 sky130_fd_sc_hd__and3_1 _2333_ (.A(net284),
    .B(net246),
    .C(\dataMemory[27][19] ),
    .X(_1493_));
 sky130_fd_sc_hd__a221o_1 _2334_ (.A1(\dataMemory[24][19] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[25][19] ),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__a211o_1 _2335_ (.A1(\dataMemory[26][19] ),
    .A2(net156),
    .B1(_1494_),
    .C1(net214),
    .X(_1495_));
 sky130_fd_sc_hd__mux4_1 _2336_ (.A0(\dataMemory[28][19] ),
    .A1(\dataMemory[29][19] ),
    .A2(\dataMemory[30][19] ),
    .A3(\dataMemory[31][19] ),
    .S0(net284),
    .S1(net246),
    .X(_1496_));
 sky130_fd_sc_hd__and3_1 _2337_ (.A(net284),
    .B(net246),
    .C(\dataMemory[7][19] ),
    .X(_1497_));
 sky130_fd_sc_hd__a221o_1 _2338_ (.A1(\dataMemory[6][19] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[5][19] ),
    .C1(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__a211o_1 _2339_ (.A1(\dataMemory[4][19] ),
    .A2(net172),
    .B1(_1498_),
    .C1(net190),
    .X(_1499_));
 sky130_fd_sc_hd__and3_1 _2340_ (.A(net285),
    .B(net247),
    .C(\dataMemory[3][19] ),
    .X(_1500_));
 sky130_fd_sc_hd__a221o_1 _2341_ (.A1(\dataMemory[2][19] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[1][19] ),
    .C1(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__a211o_1 _2342_ (.A1(\dataMemory[0][19] ),
    .A2(net172),
    .B1(_1501_),
    .C1(net214),
    .X(_1502_));
 sky130_fd_sc_hd__and3_1 _2343_ (.A(net284),
    .B(net246),
    .C(\dataMemory[11][19] ),
    .X(_1503_));
 sky130_fd_sc_hd__a221o_1 _2344_ (.A1(\dataMemory[8][19] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[9][19] ),
    .C1(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__a211o_1 _2345_ (.A1(\dataMemory[10][19] ),
    .A2(net156),
    .B1(_1504_),
    .C1(net214),
    .X(_1505_));
 sky130_fd_sc_hd__mux4_1 _2346_ (.A0(\dataMemory[12][19] ),
    .A1(\dataMemory[13][19] ),
    .A2(\dataMemory[14][19] ),
    .A3(\dataMemory[15][19] ),
    .S0(net284),
    .S1(net246),
    .X(_1506_));
 sky130_fd_sc_hd__o21a_1 _2347_ (.A1(net190),
    .A2(_1506_),
    .B1(net207),
    .X(_1507_));
 sky130_fd_sc_hd__a32o_1 _2348_ (.A1(net184),
    .A2(_1499_),
    .A3(_1502_),
    .B1(_1505_),
    .B2(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__o21a_1 _2349_ (.A1(net190),
    .A2(_1496_),
    .B1(net207),
    .X(_1509_));
 sky130_fd_sc_hd__a32o_1 _2350_ (.A1(net184),
    .A2(_1489_),
    .A3(_1492_),
    .B1(_1495_),
    .B2(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__mux2_4 _2351_ (.A0(_1508_),
    .A1(_1510_),
    .S(net203),
    .X(net50));
 sky130_fd_sc_hd__and3_1 _2352_ (.A(net285),
    .B(net247),
    .C(\dataMemory[23][20] ),
    .X(_1511_));
 sky130_fd_sc_hd__a221o_1 _2353_ (.A1(\dataMemory[22][20] ),
    .A2(net156),
    .B1(net142),
    .B2(\dataMemory[21][20] ),
    .C1(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__a211o_1 _2354_ (.A1(\dataMemory[20][20] ),
    .A2(net172),
    .B1(_1512_),
    .C1(net190),
    .X(_1513_));
 sky130_fd_sc_hd__and3_1 _2355_ (.A(net285),
    .B(net247),
    .C(\dataMemory[19][20] ),
    .X(_1514_));
 sky130_fd_sc_hd__a221o_1 _2356_ (.A1(\dataMemory[18][20] ),
    .A2(net156),
    .B1(net142),
    .B2(\dataMemory[17][20] ),
    .C1(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__a211o_1 _2357_ (.A1(\dataMemory[16][20] ),
    .A2(net172),
    .B1(_1515_),
    .C1(net214),
    .X(_1516_));
 sky130_fd_sc_hd__and3_1 _2358_ (.A(net285),
    .B(net247),
    .C(\dataMemory[27][20] ),
    .X(_1517_));
 sky130_fd_sc_hd__a221o_1 _2359_ (.A1(\dataMemory[24][20] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[25][20] ),
    .C1(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__a211o_1 _2360_ (.A1(\dataMemory[26][20] ),
    .A2(net156),
    .B1(_1518_),
    .C1(net214),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_1 _2361_ (.A0(\dataMemory[28][20] ),
    .A1(\dataMemory[29][20] ),
    .A2(\dataMemory[30][20] ),
    .A3(\dataMemory[31][20] ),
    .S0(net285),
    .S1(net247),
    .X(_1520_));
 sky130_fd_sc_hd__and3_1 _2362_ (.A(net285),
    .B(net247),
    .C(\dataMemory[7][20] ),
    .X(_1521_));
 sky130_fd_sc_hd__a221o_1 _2363_ (.A1(\dataMemory[6][20] ),
    .A2(net157),
    .B1(net142),
    .B2(\dataMemory[5][20] ),
    .C1(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__a211o_1 _2364_ (.A1(\dataMemory[4][20] ),
    .A2(net173),
    .B1(_1522_),
    .C1(net190),
    .X(_1523_));
 sky130_fd_sc_hd__and3_1 _2365_ (.A(net285),
    .B(net247),
    .C(\dataMemory[3][20] ),
    .X(_1524_));
 sky130_fd_sc_hd__a221o_1 _2366_ (.A1(\dataMemory[2][20] ),
    .A2(net157),
    .B1(net142),
    .B2(\dataMemory[1][20] ),
    .C1(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__a211o_1 _2367_ (.A1(\dataMemory[0][20] ),
    .A2(net173),
    .B1(_1525_),
    .C1(net214),
    .X(_1526_));
 sky130_fd_sc_hd__and3_1 _2368_ (.A(net285),
    .B(net247),
    .C(\dataMemory[11][20] ),
    .X(_1527_));
 sky130_fd_sc_hd__a221o_1 _2369_ (.A1(\dataMemory[8][20] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[9][20] ),
    .C1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__a211o_1 _2370_ (.A1(\dataMemory[10][20] ),
    .A2(net157),
    .B1(_1528_),
    .C1(net214),
    .X(_1529_));
 sky130_fd_sc_hd__mux4_1 _2371_ (.A0(\dataMemory[12][20] ),
    .A1(\dataMemory[13][20] ),
    .A2(\dataMemory[14][20] ),
    .A3(\dataMemory[15][20] ),
    .S0(net285),
    .S1(net247),
    .X(_1530_));
 sky130_fd_sc_hd__o21a_1 _2372_ (.A1(net190),
    .A2(_1530_),
    .B1(net207),
    .X(_1531_));
 sky130_fd_sc_hd__a32o_1 _2373_ (.A1(net184),
    .A2(_1523_),
    .A3(_1526_),
    .B1(_1529_),
    .B2(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__o21a_1 _2374_ (.A1(net190),
    .A2(_1520_),
    .B1(net207),
    .X(_1533_));
 sky130_fd_sc_hd__a32o_1 _2375_ (.A1(net184),
    .A2(_1513_),
    .A3(_1516_),
    .B1(_1519_),
    .B2(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_4 _2376_ (.A0(_1532_),
    .A1(_1534_),
    .S(net203),
    .X(net52));
 sky130_fd_sc_hd__and3_1 _2377_ (.A(net291),
    .B(net253),
    .C(\dataMemory[23][21] ),
    .X(_1535_));
 sky130_fd_sc_hd__a221o_1 _2378_ (.A1(\dataMemory[22][21] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[21][21] ),
    .C1(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__a211o_1 _2379_ (.A1(\dataMemory[20][21] ),
    .A2(net180),
    .B1(_1536_),
    .C1(net194),
    .X(_1537_));
 sky130_fd_sc_hd__and3_1 _2380_ (.A(net289),
    .B(net251),
    .C(\dataMemory[19][21] ),
    .X(_1538_));
 sky130_fd_sc_hd__a221o_1 _2381_ (.A1(\dataMemory[18][21] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[17][21] ),
    .C1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__a211o_1 _2382_ (.A1(\dataMemory[16][21] ),
    .A2(net176),
    .B1(_1539_),
    .C1(net217),
    .X(_1540_));
 sky130_fd_sc_hd__and3_1 _2383_ (.A(net288),
    .B(net251),
    .C(\dataMemory[27][21] ),
    .X(_1541_));
 sky130_fd_sc_hd__a221o_1 _2384_ (.A1(\dataMemory[24][21] ),
    .A2(net175),
    .B1(net144),
    .B2(\dataMemory[25][21] ),
    .C1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__a211o_1 _2385_ (.A1(\dataMemory[26][21] ),
    .A2(net160),
    .B1(_1542_),
    .C1(net216),
    .X(_1543_));
 sky130_fd_sc_hd__mux4_1 _2386_ (.A0(\dataMemory[28][21] ),
    .A1(\dataMemory[29][21] ),
    .A2(\dataMemory[30][21] ),
    .A3(\dataMemory[31][21] ),
    .S0(net290),
    .S1(net251),
    .X(_1544_));
 sky130_fd_sc_hd__and3_1 _2387_ (.A(net291),
    .B(net253),
    .C(\dataMemory[7][21] ),
    .X(_1545_));
 sky130_fd_sc_hd__a221o_1 _2388_ (.A1(\dataMemory[6][21] ),
    .A2(net159),
    .B1(net143),
    .B2(\dataMemory[5][21] ),
    .C1(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__a211o_1 _2389_ (.A1(\dataMemory[4][21] ),
    .A2(net175),
    .B1(_1546_),
    .C1(net191),
    .X(_1547_));
 sky130_fd_sc_hd__and3_1 _2390_ (.A(net288),
    .B(net250),
    .C(\dataMemory[3][21] ),
    .X(_1548_));
 sky130_fd_sc_hd__a221o_1 _2391_ (.A1(\dataMemory[2][21] ),
    .A2(net158),
    .B1(net143),
    .B2(\dataMemory[1][21] ),
    .C1(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__a211o_1 _2392_ (.A1(\dataMemory[0][21] ),
    .A2(net174),
    .B1(_1549_),
    .C1(net216),
    .X(_1550_));
 sky130_fd_sc_hd__and3_1 _2393_ (.A(net2),
    .B(net250),
    .C(\dataMemory[11][21] ),
    .X(_1551_));
 sky130_fd_sc_hd__a221o_1 _2394_ (.A1(\dataMemory[8][21] ),
    .A2(net174),
    .B1(net143),
    .B2(\dataMemory[9][21] ),
    .C1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__a211o_1 _2395_ (.A1(\dataMemory[10][21] ),
    .A2(net158),
    .B1(_1552_),
    .C1(net216),
    .X(_1553_));
 sky130_fd_sc_hd__mux4_1 _2396_ (.A0(\dataMemory[12][21] ),
    .A1(\dataMemory[13][21] ),
    .A2(\dataMemory[14][21] ),
    .A3(\dataMemory[15][21] ),
    .S0(net2),
    .S1(net250),
    .X(_1554_));
 sky130_fd_sc_hd__o21a_1 _2397_ (.A1(net191),
    .A2(_1554_),
    .B1(net209),
    .X(_1555_));
 sky130_fd_sc_hd__a32o_1 _2398_ (.A1(net186),
    .A2(_1547_),
    .A3(_1550_),
    .B1(_1553_),
    .B2(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__o21a_1 _2399_ (.A1(net192),
    .A2(_1544_),
    .B1(net209),
    .X(_1557_));
 sky130_fd_sc_hd__a32o_1 _2400_ (.A1(net186),
    .A2(_1537_),
    .A3(_1540_),
    .B1(_1543_),
    .B2(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_2 _2401_ (.A0(_1556_),
    .A1(_1558_),
    .S(net204),
    .X(net53));
 sky130_fd_sc_hd__and3_1 _2402_ (.A(net291),
    .B(net253),
    .C(\dataMemory[23][22] ),
    .X(_1559_));
 sky130_fd_sc_hd__a221o_1 _2403_ (.A1(\dataMemory[22][22] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[21][22] ),
    .C1(_1559_),
    .X(_1560_));
 sky130_fd_sc_hd__a211o_1 _2404_ (.A1(\dataMemory[20][22] ),
    .A2(net179),
    .B1(_1560_),
    .C1(net193),
    .X(_1561_));
 sky130_fd_sc_hd__and3_1 _2405_ (.A(net291),
    .B(net253),
    .C(\dataMemory[19][22] ),
    .X(_1562_));
 sky130_fd_sc_hd__a221o_1 _2406_ (.A1(\dataMemory[18][22] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[17][22] ),
    .C1(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a211o_1 _2407_ (.A1(\dataMemory[16][22] ),
    .A2(net179),
    .B1(_1563_),
    .C1(net218),
    .X(_1564_));
 sky130_fd_sc_hd__and3_1 _2408_ (.A(net291),
    .B(net253),
    .C(\dataMemory[27][22] ),
    .X(_1565_));
 sky130_fd_sc_hd__a221o_1 _2409_ (.A1(\dataMemory[24][22] ),
    .A2(net179),
    .B1(net146),
    .B2(\dataMemory[25][22] ),
    .C1(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__a211o_1 _2410_ (.A1(\dataMemory[26][22] ),
    .A2(net162),
    .B1(_1566_),
    .C1(net218),
    .X(_1567_));
 sky130_fd_sc_hd__mux4_1 _2411_ (.A0(\dataMemory[28][22] ),
    .A1(\dataMemory[29][22] ),
    .A2(\dataMemory[30][22] ),
    .A3(\dataMemory[31][22] ),
    .S0(net291),
    .S1(net253),
    .X(_1568_));
 sky130_fd_sc_hd__and3_1 _2412_ (.A(net292),
    .B(net254),
    .C(\dataMemory[7][22] ),
    .X(_1569_));
 sky130_fd_sc_hd__a221o_1 _2413_ (.A1(\dataMemory[6][22] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[5][22] ),
    .C1(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__a211o_1 _2414_ (.A1(\dataMemory[4][22] ),
    .A2(net178),
    .B1(_1570_),
    .C1(net193),
    .X(_1571_));
 sky130_fd_sc_hd__and3_1 _2415_ (.A(net292),
    .B(net254),
    .C(\dataMemory[3][22] ),
    .X(_1572_));
 sky130_fd_sc_hd__a221o_1 _2416_ (.A1(\dataMemory[2][22] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[1][22] ),
    .C1(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__a211o_1 _2417_ (.A1(\dataMemory[0][22] ),
    .A2(net178),
    .B1(_1573_),
    .C1(net219),
    .X(_1574_));
 sky130_fd_sc_hd__and3_1 _2418_ (.A(net292),
    .B(net254),
    .C(\dataMemory[11][22] ),
    .X(_1575_));
 sky130_fd_sc_hd__a221o_1 _2419_ (.A1(\dataMemory[8][22] ),
    .A2(net178),
    .B1(net147),
    .B2(\dataMemory[9][22] ),
    .C1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__a211o_1 _2420_ (.A1(\dataMemory[10][22] ),
    .A2(net163),
    .B1(_1576_),
    .C1(net219),
    .X(_1577_));
 sky130_fd_sc_hd__mux4_1 _2421_ (.A0(\dataMemory[12][22] ),
    .A1(\dataMemory[13][22] ),
    .A2(\dataMemory[14][22] ),
    .A3(\dataMemory[15][22] ),
    .S0(net292),
    .S1(net254),
    .X(_1578_));
 sky130_fd_sc_hd__o21a_1 _2422_ (.A1(net193),
    .A2(_1578_),
    .B1(net208),
    .X(_1579_));
 sky130_fd_sc_hd__a32o_1 _2423_ (.A1(net185),
    .A2(_1571_),
    .A3(_1574_),
    .B1(_1577_),
    .B2(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__o21a_1 _2424_ (.A1(net193),
    .A2(_1568_),
    .B1(net208),
    .X(_1581_));
 sky130_fd_sc_hd__a32o_1 _2425_ (.A1(net185),
    .A2(_1561_),
    .A3(_1564_),
    .B1(_1567_),
    .B2(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_2 _2426_ (.A0(_1580_),
    .A1(_1582_),
    .S(net204),
    .X(net54));
 sky130_fd_sc_hd__and3_1 _2427_ (.A(net291),
    .B(net253),
    .C(\dataMemory[23][23] ),
    .X(_1583_));
 sky130_fd_sc_hd__a221o_1 _2428_ (.A1(\dataMemory[22][23] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[21][23] ),
    .C1(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__a211o_1 _2429_ (.A1(\dataMemory[20][23] ),
    .A2(net179),
    .B1(_1584_),
    .C1(net193),
    .X(_1585_));
 sky130_fd_sc_hd__and3_1 _2430_ (.A(net291),
    .B(net253),
    .C(\dataMemory[19][23] ),
    .X(_1586_));
 sky130_fd_sc_hd__a221o_1 _2431_ (.A1(\dataMemory[18][23] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[17][23] ),
    .C1(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__a211o_1 _2432_ (.A1(\dataMemory[16][23] ),
    .A2(net179),
    .B1(_1587_),
    .C1(net219),
    .X(_1588_));
 sky130_fd_sc_hd__and3_1 _2433_ (.A(net291),
    .B(net253),
    .C(\dataMemory[27][23] ),
    .X(_1589_));
 sky130_fd_sc_hd__a221o_1 _2434_ (.A1(\dataMemory[24][23] ),
    .A2(net179),
    .B1(net146),
    .B2(\dataMemory[25][23] ),
    .C1(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__a211o_1 _2435_ (.A1(\dataMemory[26][23] ),
    .A2(net162),
    .B1(_1590_),
    .C1(net218),
    .X(_1591_));
 sky130_fd_sc_hd__mux4_1 _2436_ (.A0(\dataMemory[28][23] ),
    .A1(\dataMemory[29][23] ),
    .A2(\dataMemory[30][23] ),
    .A3(\dataMemory[31][23] ),
    .S0(net291),
    .S1(net253),
    .X(_1592_));
 sky130_fd_sc_hd__and3_1 _2437_ (.A(net292),
    .B(net254),
    .C(\dataMemory[7][23] ),
    .X(_1593_));
 sky130_fd_sc_hd__a221o_1 _2438_ (.A1(\dataMemory[6][23] ),
    .A2(net163),
    .B1(net147),
    .B2(\dataMemory[5][23] ),
    .C1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__a211o_1 _2439_ (.A1(\dataMemory[4][23] ),
    .A2(net178),
    .B1(_1594_),
    .C1(net193),
    .X(_1595_));
 sky130_fd_sc_hd__and3_1 _2440_ (.A(net292),
    .B(net254),
    .C(\dataMemory[3][23] ),
    .X(_1596_));
 sky130_fd_sc_hd__a221o_1 _2441_ (.A1(\dataMemory[2][23] ),
    .A2(net162),
    .B1(net147),
    .B2(\dataMemory[1][23] ),
    .C1(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__a211o_1 _2442_ (.A1(\dataMemory[0][23] ),
    .A2(net178),
    .B1(_1597_),
    .C1(net219),
    .X(_1598_));
 sky130_fd_sc_hd__and3_1 _2443_ (.A(net292),
    .B(net254),
    .C(\dataMemory[11][23] ),
    .X(_1599_));
 sky130_fd_sc_hd__a221o_1 _2444_ (.A1(\dataMemory[8][23] ),
    .A2(net178),
    .B1(net146),
    .B2(\dataMemory[9][23] ),
    .C1(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__a211o_1 _2445_ (.A1(\dataMemory[10][23] ),
    .A2(net162),
    .B1(_1600_),
    .C1(net219),
    .X(_1601_));
 sky130_fd_sc_hd__mux4_1 _2446_ (.A0(\dataMemory[12][23] ),
    .A1(\dataMemory[13][23] ),
    .A2(\dataMemory[14][23] ),
    .A3(\dataMemory[15][23] ),
    .S0(net292),
    .S1(net254),
    .X(_1602_));
 sky130_fd_sc_hd__o21a_1 _2447_ (.A1(net193),
    .A2(_1602_),
    .B1(net208),
    .X(_1603_));
 sky130_fd_sc_hd__a32o_1 _2448_ (.A1(net185),
    .A2(_1595_),
    .A3(_1598_),
    .B1(_1601_),
    .B2(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__o21a_1 _2449_ (.A1(net193),
    .A2(_1592_),
    .B1(net208),
    .X(_1605_));
 sky130_fd_sc_hd__a32o_1 _2450_ (.A1(net185),
    .A2(_1585_),
    .A3(_1588_),
    .B1(_1591_),
    .B2(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__mux2_2 _2451_ (.A0(_1604_),
    .A1(_1606_),
    .S(net204),
    .X(net55));
 sky130_fd_sc_hd__and3_1 _2452_ (.A(net291),
    .B(net253),
    .C(\dataMemory[23][24] ),
    .X(_1607_));
 sky130_fd_sc_hd__a221o_1 _2453_ (.A1(\dataMemory[22][24] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[21][24] ),
    .C1(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__a211o_1 _2454_ (.A1(\dataMemory[20][24] ),
    .A2(net179),
    .B1(_1608_),
    .C1(net193),
    .X(_1609_));
 sky130_fd_sc_hd__and3_1 _2455_ (.A(net295),
    .B(net257),
    .C(\dataMemory[19][24] ),
    .X(_1610_));
 sky130_fd_sc_hd__a221o_1 _2456_ (.A1(\dataMemory[18][24] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[17][24] ),
    .C1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__a211o_1 _2457_ (.A1(\dataMemory[16][24] ),
    .A2(net180),
    .B1(_1611_),
    .C1(net220),
    .X(_1612_));
 sky130_fd_sc_hd__and3_1 _2458_ (.A(net295),
    .B(net257),
    .C(\dataMemory[27][24] ),
    .X(_1613_));
 sky130_fd_sc_hd__a221o_1 _2459_ (.A1(\dataMemory[24][24] ),
    .A2(net179),
    .B1(net146),
    .B2(\dataMemory[25][24] ),
    .C1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__a211o_1 _2460_ (.A1(\dataMemory[26][24] ),
    .A2(net162),
    .B1(_1614_),
    .C1(net218),
    .X(_1615_));
 sky130_fd_sc_hd__mux4_1 _2461_ (.A0(\dataMemory[28][24] ),
    .A1(\dataMemory[29][24] ),
    .A2(\dataMemory[30][24] ),
    .A3(\dataMemory[31][24] ),
    .S0(net294),
    .S1(net256),
    .X(_1616_));
 sky130_fd_sc_hd__and3_1 _2462_ (.A(net292),
    .B(net254),
    .C(\dataMemory[7][24] ),
    .X(_1617_));
 sky130_fd_sc_hd__a221o_1 _2463_ (.A1(\dataMemory[6][24] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[5][24] ),
    .C1(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__a211o_1 _2464_ (.A1(\dataMemory[4][24] ),
    .A2(net178),
    .B1(_1618_),
    .C1(net193),
    .X(_1619_));
 sky130_fd_sc_hd__and3_1 _2465_ (.A(net292),
    .B(net254),
    .C(\dataMemory[3][24] ),
    .X(_1620_));
 sky130_fd_sc_hd__a221o_1 _2466_ (.A1(\dataMemory[2][24] ),
    .A2(net162),
    .B1(net146),
    .B2(\dataMemory[1][24] ),
    .C1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__a211o_1 _2467_ (.A1(\dataMemory[0][24] ),
    .A2(net178),
    .B1(_1621_),
    .C1(net219),
    .X(_1622_));
 sky130_fd_sc_hd__and3_1 _2468_ (.A(net295),
    .B(net257),
    .C(\dataMemory[11][24] ),
    .X(_1623_));
 sky130_fd_sc_hd__a221o_1 _2469_ (.A1(\dataMemory[8][24] ),
    .A2(net178),
    .B1(net146),
    .B2(\dataMemory[9][24] ),
    .C1(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__a211o_1 _2470_ (.A1(\dataMemory[10][24] ),
    .A2(net162),
    .B1(_1624_),
    .C1(net219),
    .X(_1625_));
 sky130_fd_sc_hd__mux4_1 _2471_ (.A0(\dataMemory[12][24] ),
    .A1(\dataMemory[13][24] ),
    .A2(\dataMemory[14][24] ),
    .A3(\dataMemory[15][24] ),
    .S0(net295),
    .S1(net257),
    .X(_1626_));
 sky130_fd_sc_hd__o21a_1 _2472_ (.A1(net193),
    .A2(_1626_),
    .B1(net208),
    .X(_1627_));
 sky130_fd_sc_hd__a32o_1 _2473_ (.A1(net185),
    .A2(_1619_),
    .A3(_1622_),
    .B1(_1625_),
    .B2(_1627_),
    .X(_1628_));
 sky130_fd_sc_hd__o21a_1 _2474_ (.A1(net194),
    .A2(_1616_),
    .B1(net208),
    .X(_1629_));
 sky130_fd_sc_hd__a32o_1 _2475_ (.A1(net185),
    .A2(_1609_),
    .A3(_1612_),
    .B1(_1615_),
    .B2(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_2 _2476_ (.A0(_1628_),
    .A1(_1630_),
    .S(net204),
    .X(net56));
 sky130_fd_sc_hd__and3_1 _2477_ (.A(net290),
    .B(net251),
    .C(\dataMemory[23][25] ),
    .X(_1631_));
 sky130_fd_sc_hd__a221o_1 _2478_ (.A1(\dataMemory[22][25] ),
    .A2(net161),
    .B1(net145),
    .B2(\dataMemory[21][25] ),
    .C1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__a211o_1 _2479_ (.A1(\dataMemory[20][25] ),
    .A2(net177),
    .B1(_1632_),
    .C1(net192),
    .X(_1633_));
 sky130_fd_sc_hd__and3_1 _2480_ (.A(net290),
    .B(net251),
    .C(\dataMemory[19][25] ),
    .X(_1634_));
 sky130_fd_sc_hd__a221o_1 _2481_ (.A1(\dataMemory[18][25] ),
    .A2(net161),
    .B1(net145),
    .B2(\dataMemory[17][25] ),
    .C1(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__a211o_1 _2482_ (.A1(\dataMemory[16][25] ),
    .A2(net177),
    .B1(_1635_),
    .C1(net217),
    .X(_1636_));
 sky130_fd_sc_hd__and3_1 _2483_ (.A(net290),
    .B(net251),
    .C(\dataMemory[27][25] ),
    .X(_1637_));
 sky130_fd_sc_hd__a221o_1 _2484_ (.A1(\dataMemory[24][25] ),
    .A2(net177),
    .B1(net145),
    .B2(\dataMemory[25][25] ),
    .C1(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__a211o_1 _2485_ (.A1(\dataMemory[26][25] ),
    .A2(net161),
    .B1(_1638_),
    .C1(net217),
    .X(_1639_));
 sky130_fd_sc_hd__mux4_1 _2486_ (.A0(\dataMemory[28][25] ),
    .A1(\dataMemory[29][25] ),
    .A2(\dataMemory[30][25] ),
    .A3(\dataMemory[31][25] ),
    .S0(net290),
    .S1(net251),
    .X(_1640_));
 sky130_fd_sc_hd__and3_1 _2487_ (.A(net290),
    .B(net251),
    .C(\dataMemory[7][25] ),
    .X(_1641_));
 sky130_fd_sc_hd__a221o_1 _2488_ (.A1(\dataMemory[6][25] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[5][25] ),
    .C1(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__a211o_1 _2489_ (.A1(\dataMemory[4][25] ),
    .A2(net176),
    .B1(_1642_),
    .C1(net192),
    .X(_1643_));
 sky130_fd_sc_hd__and3_1 _2490_ (.A(net290),
    .B(net251),
    .C(\dataMemory[3][25] ),
    .X(_1644_));
 sky130_fd_sc_hd__a221o_1 _2491_ (.A1(\dataMemory[2][25] ),
    .A2(net161),
    .B1(net144),
    .B2(\dataMemory[1][25] ),
    .C1(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__a211o_1 _2492_ (.A1(\dataMemory[0][25] ),
    .A2(net180),
    .B1(_1645_),
    .C1(net220),
    .X(_1646_));
 sky130_fd_sc_hd__and3_1 _2493_ (.A(net290),
    .B(net251),
    .C(\dataMemory[11][25] ),
    .X(_1647_));
 sky130_fd_sc_hd__a221o_1 _2494_ (.A1(\dataMemory[8][25] ),
    .A2(net176),
    .B1(net144),
    .B2(\dataMemory[9][25] ),
    .C1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__a211o_1 _2495_ (.A1(\dataMemory[10][25] ),
    .A2(net160),
    .B1(_1648_),
    .C1(net217),
    .X(_1649_));
 sky130_fd_sc_hd__mux4_1 _2496_ (.A0(\dataMemory[12][25] ),
    .A1(\dataMemory[13][25] ),
    .A2(\dataMemory[14][25] ),
    .A3(\dataMemory[15][25] ),
    .S0(net290),
    .S1(net251),
    .X(_1650_));
 sky130_fd_sc_hd__o21a_1 _2497_ (.A1(net192),
    .A2(_1650_),
    .B1(net208),
    .X(_1651_));
 sky130_fd_sc_hd__a32o_1 _2498_ (.A1(net186),
    .A2(_1643_),
    .A3(_1646_),
    .B1(_1649_),
    .B2(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__o21a_1 _2499_ (.A1(net192),
    .A2(_1640_),
    .B1(net208),
    .X(_1653_));
 sky130_fd_sc_hd__a32o_1 _2500_ (.A1(net186),
    .A2(_1633_),
    .A3(_1636_),
    .B1(_1639_),
    .B2(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__mux2_2 _2501_ (.A0(_1652_),
    .A1(_1654_),
    .S(net204),
    .X(net57));
 sky130_fd_sc_hd__and3_1 _2502_ (.A(net285),
    .B(net247),
    .C(\dataMemory[23][26] ),
    .X(_1655_));
 sky130_fd_sc_hd__a221o_1 _2503_ (.A1(\dataMemory[22][26] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[21][26] ),
    .C1(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__a211o_1 _2504_ (.A1(\dataMemory[20][26] ),
    .A2(net172),
    .B1(_1656_),
    .C1(net190),
    .X(_1657_));
 sky130_fd_sc_hd__and3_1 _2505_ (.A(net289),
    .B(net252),
    .C(\dataMemory[19][26] ),
    .X(_1658_));
 sky130_fd_sc_hd__a221o_1 _2506_ (.A1(\dataMemory[18][26] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[17][26] ),
    .C1(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__a211o_1 _2507_ (.A1(\dataMemory[16][26] ),
    .A2(net176),
    .B1(_1659_),
    .C1(net217),
    .X(_1660_));
 sky130_fd_sc_hd__and3_1 _2508_ (.A(net285),
    .B(net247),
    .C(\dataMemory[27][26] ),
    .X(_1661_));
 sky130_fd_sc_hd__a221o_1 _2509_ (.A1(\dataMemory[24][26] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[25][26] ),
    .C1(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__a211o_1 _2510_ (.A1(\dataMemory[26][26] ),
    .A2(net157),
    .B1(_1662_),
    .C1(net214),
    .X(_1663_));
 sky130_fd_sc_hd__mux4_1 _2511_ (.A0(\dataMemory[28][26] ),
    .A1(\dataMemory[29][26] ),
    .A2(\dataMemory[30][26] ),
    .A3(\dataMemory[31][26] ),
    .S0(net285),
    .S1(net247),
    .X(_1664_));
 sky130_fd_sc_hd__and3_1 _2512_ (.A(net289),
    .B(net252),
    .C(\dataMemory[7][26] ),
    .X(_1665_));
 sky130_fd_sc_hd__a221o_1 _2513_ (.A1(\dataMemory[6][26] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[5][26] ),
    .C1(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__a211o_1 _2514_ (.A1(\dataMemory[4][26] ),
    .A2(net176),
    .B1(_1666_),
    .C1(net189),
    .X(_1667_));
 sky130_fd_sc_hd__and3_1 _2515_ (.A(net289),
    .B(net252),
    .C(\dataMemory[3][26] ),
    .X(_1668_));
 sky130_fd_sc_hd__a221o_1 _2516_ (.A1(\dataMemory[2][26] ),
    .A2(net156),
    .B1(net141),
    .B2(\dataMemory[1][26] ),
    .C1(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__a211o_1 _2517_ (.A1(\dataMemory[0][26] ),
    .A2(net176),
    .B1(_1669_),
    .C1(net217),
    .X(_1670_));
 sky130_fd_sc_hd__and3_1 _2518_ (.A(net286),
    .B(net248),
    .C(\dataMemory[11][26] ),
    .X(_1671_));
 sky130_fd_sc_hd__a221o_1 _2519_ (.A1(\dataMemory[8][26] ),
    .A2(net172),
    .B1(net141),
    .B2(\dataMemory[9][26] ),
    .C1(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__a211o_1 _2520_ (.A1(\dataMemory[10][26] ),
    .A2(net156),
    .B1(_1672_),
    .C1(net214),
    .X(_1673_));
 sky130_fd_sc_hd__mux4_1 _2521_ (.A0(\dataMemory[12][26] ),
    .A1(\dataMemory[13][26] ),
    .A2(\dataMemory[14][26] ),
    .A3(\dataMemory[15][26] ),
    .S0(net286),
    .S1(net248),
    .X(_1674_));
 sky130_fd_sc_hd__o21a_1 _2522_ (.A1(net189),
    .A2(_1674_),
    .B1(net209),
    .X(_1675_));
 sky130_fd_sc_hd__a32o_1 _2523_ (.A1(net184),
    .A2(_1667_),
    .A3(_1670_),
    .B1(_1673_),
    .B2(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__o21a_1 _2524_ (.A1(net190),
    .A2(_1664_),
    .B1(net209),
    .X(_1677_));
 sky130_fd_sc_hd__a32o_1 _2525_ (.A1(net184),
    .A2(_1657_),
    .A3(_1660_),
    .B1(_1663_),
    .B2(_1677_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_4 _2526_ (.A0(_1676_),
    .A1(_1678_),
    .S(net205),
    .X(net58));
 sky130_fd_sc_hd__and3_1 _2527_ (.A(net290),
    .B(net251),
    .C(\dataMemory[23][27] ),
    .X(_1679_));
 sky130_fd_sc_hd__a221o_1 _2528_ (.A1(\dataMemory[22][27] ),
    .A2(net160),
    .B1(net144),
    .B2(\dataMemory[21][27] ),
    .C1(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__a211o_1 _2529_ (.A1(\dataMemory[20][27] ),
    .A2(net177),
    .B1(_1680_),
    .C1(net192),
    .X(_1681_));
 sky130_fd_sc_hd__and3_1 _2530_ (.A(net290),
    .B(net251),
    .C(\dataMemory[19][27] ),
    .X(_1682_));
 sky130_fd_sc_hd__a221o_1 _2531_ (.A1(\dataMemory[18][27] ),
    .A2(net161),
    .B1(net145),
    .B2(\dataMemory[17][27] ),
    .C1(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__a211o_1 _2532_ (.A1(\dataMemory[16][27] ),
    .A2(net176),
    .B1(_1683_),
    .C1(net217),
    .X(_1684_));
 sky130_fd_sc_hd__and3_1 _2533_ (.A(net289),
    .B(net252),
    .C(\dataMemory[27][27] ),
    .X(_1685_));
 sky130_fd_sc_hd__a221o_1 _2534_ (.A1(\dataMemory[24][27] ),
    .A2(net176),
    .B1(net144),
    .B2(\dataMemory[25][27] ),
    .C1(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__a211o_1 _2535_ (.A1(\dataMemory[26][27] ),
    .A2(net161),
    .B1(_1686_),
    .C1(net217),
    .X(_1687_));
 sky130_fd_sc_hd__mux4_1 _2536_ (.A0(\dataMemory[28][27] ),
    .A1(\dataMemory[29][27] ),
    .A2(\dataMemory[30][27] ),
    .A3(\dataMemory[31][27] ),
    .S0(net290),
    .S1(net251),
    .X(_1688_));
 sky130_fd_sc_hd__and3_1 _2537_ (.A(net290),
    .B(net251),
    .C(\dataMemory[7][27] ),
    .X(_1689_));
 sky130_fd_sc_hd__a221o_1 _2538_ (.A1(\dataMemory[6][27] ),
    .A2(net160),
    .B1(net145),
    .B2(\dataMemory[5][27] ),
    .C1(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__a211o_1 _2539_ (.A1(\dataMemory[4][27] ),
    .A2(net176),
    .B1(_1690_),
    .C1(net192),
    .X(_1691_));
 sky130_fd_sc_hd__and3_1 _2540_ (.A(net290),
    .B(net3),
    .C(\dataMemory[3][27] ),
    .X(_1692_));
 sky130_fd_sc_hd__a221o_1 _2541_ (.A1(\dataMemory[2][27] ),
    .A2(net160),
    .B1(net145),
    .B2(\dataMemory[1][27] ),
    .C1(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__a211o_1 _2542_ (.A1(\dataMemory[0][27] ),
    .A2(net177),
    .B1(_1693_),
    .C1(net217),
    .X(_1694_));
 sky130_fd_sc_hd__and3_1 _2543_ (.A(net289),
    .B(net252),
    .C(\dataMemory[11][27] ),
    .X(_1695_));
 sky130_fd_sc_hd__a221o_1 _2544_ (.A1(\dataMemory[8][27] ),
    .A2(net177),
    .B1(net144),
    .B2(\dataMemory[9][27] ),
    .C1(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__a211o_1 _2545_ (.A1(\dataMemory[10][27] ),
    .A2(net160),
    .B1(_1696_),
    .C1(net217),
    .X(_1697_));
 sky130_fd_sc_hd__mux4_1 _2546_ (.A0(\dataMemory[12][27] ),
    .A1(\dataMemory[13][27] ),
    .A2(\dataMemory[14][27] ),
    .A3(\dataMemory[15][27] ),
    .S0(net290),
    .S1(net251),
    .X(_1698_));
 sky130_fd_sc_hd__o21a_1 _2547_ (.A1(net192),
    .A2(_1698_),
    .B1(net209),
    .X(_1699_));
 sky130_fd_sc_hd__a32o_1 _2548_ (.A1(net186),
    .A2(_1691_),
    .A3(_1694_),
    .B1(_1697_),
    .B2(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__o21a_1 _2549_ (.A1(net192),
    .A2(_1688_),
    .B1(net209),
    .X(_1701_));
 sky130_fd_sc_hd__a32o_1 _2550_ (.A1(net186),
    .A2(_1681_),
    .A3(_1684_),
    .B1(_1687_),
    .B2(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__mux2_2 _2551_ (.A0(_1700_),
    .A1(_1702_),
    .S(net204),
    .X(net59));
 sky130_fd_sc_hd__and3_1 _2552_ (.A(net294),
    .B(net256),
    .C(\dataMemory[23][28] ),
    .X(_1703_));
 sky130_fd_sc_hd__a221o_1 _2553_ (.A1(\dataMemory[22][28] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[21][28] ),
    .C1(_1703_),
    .X(_1704_));
 sky130_fd_sc_hd__a211o_1 _2554_ (.A1(\dataMemory[20][28] ),
    .A2(net180),
    .B1(_1704_),
    .C1(net194),
    .X(_1705_));
 sky130_fd_sc_hd__and3_1 _2555_ (.A(net294),
    .B(net256),
    .C(\dataMemory[19][28] ),
    .X(_1706_));
 sky130_fd_sc_hd__a221o_1 _2556_ (.A1(\dataMemory[18][28] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[17][28] ),
    .C1(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__a211o_1 _2557_ (.A1(\dataMemory[16][28] ),
    .A2(net180),
    .B1(_1707_),
    .C1(net220),
    .X(_1708_));
 sky130_fd_sc_hd__and3_1 _2558_ (.A(net294),
    .B(net256),
    .C(\dataMemory[27][28] ),
    .X(_1709_));
 sky130_fd_sc_hd__a221o_1 _2559_ (.A1(\dataMemory[24][28] ),
    .A2(net180),
    .B1(net148),
    .B2(\dataMemory[25][28] ),
    .C1(_1709_),
    .X(_1710_));
 sky130_fd_sc_hd__a211o_1 _2560_ (.A1(\dataMemory[26][28] ),
    .A2(net164),
    .B1(_1710_),
    .C1(net220),
    .X(_1711_));
 sky130_fd_sc_hd__mux4_1 _2561_ (.A0(\dataMemory[28][28] ),
    .A1(\dataMemory[29][28] ),
    .A2(\dataMemory[30][28] ),
    .A3(\dataMemory[31][28] ),
    .S0(net294),
    .S1(net256),
    .X(_1712_));
 sky130_fd_sc_hd__and3_1 _2562_ (.A(net294),
    .B(net256),
    .C(\dataMemory[7][28] ),
    .X(_1713_));
 sky130_fd_sc_hd__a221o_1 _2563_ (.A1(\dataMemory[6][28] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[5][28] ),
    .C1(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__a211o_1 _2564_ (.A1(\dataMemory[4][28] ),
    .A2(net180),
    .B1(_1714_),
    .C1(net194),
    .X(_1715_));
 sky130_fd_sc_hd__and3_1 _2565_ (.A(net294),
    .B(net256),
    .C(\dataMemory[3][28] ),
    .X(_1716_));
 sky130_fd_sc_hd__a221o_1 _2566_ (.A1(\dataMemory[2][28] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[1][28] ),
    .C1(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__a211o_1 _2567_ (.A1(\dataMemory[0][28] ),
    .A2(net180),
    .B1(_1717_),
    .C1(net220),
    .X(_1718_));
 sky130_fd_sc_hd__and3_1 _2568_ (.A(net294),
    .B(net256),
    .C(\dataMemory[11][28] ),
    .X(_1719_));
 sky130_fd_sc_hd__a221o_1 _2569_ (.A1(\dataMemory[8][28] ),
    .A2(net180),
    .B1(net148),
    .B2(\dataMemory[9][28] ),
    .C1(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__a211o_1 _2570_ (.A1(\dataMemory[10][28] ),
    .A2(net164),
    .B1(_1720_),
    .C1(net220),
    .X(_1721_));
 sky130_fd_sc_hd__mux4_1 _2571_ (.A0(\dataMemory[12][28] ),
    .A1(\dataMemory[13][28] ),
    .A2(\dataMemory[14][28] ),
    .A3(\dataMemory[15][28] ),
    .S0(net294),
    .S1(net256),
    .X(_1722_));
 sky130_fd_sc_hd__o21a_1 _2572_ (.A1(net194),
    .A2(_1722_),
    .B1(net208),
    .X(_1723_));
 sky130_fd_sc_hd__a32o_1 _2573_ (.A1(_1025_),
    .A2(_1715_),
    .A3(_1718_),
    .B1(_1721_),
    .B2(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__o21a_1 _2574_ (.A1(net194),
    .A2(_1712_),
    .B1(net210),
    .X(_1725_));
 sky130_fd_sc_hd__a32o_1 _2575_ (.A1(_1025_),
    .A2(_1705_),
    .A3(_1708_),
    .B1(_1711_),
    .B2(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__mux2_2 _2576_ (.A0(_1724_),
    .A1(_1726_),
    .S(net204),
    .X(net60));
 sky130_fd_sc_hd__and3_1 _2577_ (.A(net294),
    .B(net256),
    .C(\dataMemory[23][29] ),
    .X(_1727_));
 sky130_fd_sc_hd__a221o_1 _2578_ (.A1(\dataMemory[22][29] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[21][29] ),
    .C1(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__a211o_1 _2579_ (.A1(\dataMemory[20][29] ),
    .A2(net181),
    .B1(_1728_),
    .C1(net195),
    .X(_1729_));
 sky130_fd_sc_hd__and3_1 _2580_ (.A(net293),
    .B(net255),
    .C(\dataMemory[19][29] ),
    .X(_1730_));
 sky130_fd_sc_hd__a221o_1 _2581_ (.A1(\dataMemory[18][29] ),
    .A2(net165),
    .B1(net149),
    .B2(\dataMemory[17][29] ),
    .C1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__a211o_1 _2582_ (.A1(\dataMemory[16][29] ),
    .A2(net181),
    .B1(_1731_),
    .C1(net220),
    .X(_1732_));
 sky130_fd_sc_hd__and3_1 _2583_ (.A(net293),
    .B(net255),
    .C(\dataMemory[27][29] ),
    .X(_1733_));
 sky130_fd_sc_hd__a221o_1 _2584_ (.A1(\dataMemory[24][29] ),
    .A2(net181),
    .B1(net149),
    .B2(\dataMemory[25][29] ),
    .C1(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__a211o_1 _2585_ (.A1(\dataMemory[26][29] ),
    .A2(net165),
    .B1(_1734_),
    .C1(net220),
    .X(_1735_));
 sky130_fd_sc_hd__mux4_1 _2586_ (.A0(\dataMemory[28][29] ),
    .A1(\dataMemory[29][29] ),
    .A2(\dataMemory[30][29] ),
    .A3(\dataMemory[31][29] ),
    .S0(net293),
    .S1(net255),
    .X(_1736_));
 sky130_fd_sc_hd__and3_1 _2587_ (.A(net293),
    .B(net255),
    .C(\dataMemory[7][29] ),
    .X(_1737_));
 sky130_fd_sc_hd__a221o_1 _2588_ (.A1(\dataMemory[6][29] ),
    .A2(net165),
    .B1(net149),
    .B2(\dataMemory[5][29] ),
    .C1(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__a211o_1 _2589_ (.A1(\dataMemory[4][29] ),
    .A2(net181),
    .B1(_1738_),
    .C1(net195),
    .X(_1739_));
 sky130_fd_sc_hd__and3_1 _2590_ (.A(net293),
    .B(net255),
    .C(\dataMemory[3][29] ),
    .X(_1740_));
 sky130_fd_sc_hd__a221o_1 _2591_ (.A1(\dataMemory[2][29] ),
    .A2(net165),
    .B1(net149),
    .B2(\dataMemory[1][29] ),
    .C1(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__a211o_1 _2592_ (.A1(\dataMemory[0][29] ),
    .A2(net181),
    .B1(_1741_),
    .C1(net220),
    .X(_1742_));
 sky130_fd_sc_hd__and3_1 _2593_ (.A(net293),
    .B(net255),
    .C(\dataMemory[11][29] ),
    .X(_1743_));
 sky130_fd_sc_hd__a221o_1 _2594_ (.A1(\dataMemory[8][29] ),
    .A2(net181),
    .B1(net149),
    .B2(\dataMemory[9][29] ),
    .C1(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__a211o_1 _2595_ (.A1(\dataMemory[10][29] ),
    .A2(net165),
    .B1(_1744_),
    .C1(net220),
    .X(_1745_));
 sky130_fd_sc_hd__mux4_1 _2596_ (.A0(\dataMemory[12][29] ),
    .A1(\dataMemory[13][29] ),
    .A2(\dataMemory[14][29] ),
    .A3(\dataMemory[15][29] ),
    .S0(net293),
    .S1(net255),
    .X(_1746_));
 sky130_fd_sc_hd__o21a_1 _2597_ (.A1(net194),
    .A2(_1746_),
    .B1(net210),
    .X(_1747_));
 sky130_fd_sc_hd__a32o_1 _2598_ (.A1(_1025_),
    .A2(_1739_),
    .A3(_1742_),
    .B1(_1745_),
    .B2(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__o21a_1 _2599_ (.A1(net194),
    .A2(_1736_),
    .B1(net210),
    .X(_1749_));
 sky130_fd_sc_hd__a32o_1 _2600_ (.A1(net185),
    .A2(_1729_),
    .A3(_1732_),
    .B1(_1735_),
    .B2(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(_1748_),
    .A1(_1750_),
    .S(net204),
    .X(net61));
 sky130_fd_sc_hd__and3_1 _2602_ (.A(net294),
    .B(net256),
    .C(\dataMemory[23][30] ),
    .X(_1751_));
 sky130_fd_sc_hd__a221o_1 _2603_ (.A1(\dataMemory[22][30] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[21][30] ),
    .C1(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a211o_1 _2604_ (.A1(\dataMemory[20][30] ),
    .A2(net180),
    .B1(_1752_),
    .C1(net194),
    .X(_1753_));
 sky130_fd_sc_hd__and3_1 _2605_ (.A(net293),
    .B(net255),
    .C(\dataMemory[19][30] ),
    .X(_1754_));
 sky130_fd_sc_hd__a221o_1 _2606_ (.A1(\dataMemory[18][30] ),
    .A2(net165),
    .B1(net149),
    .B2(\dataMemory[17][30] ),
    .C1(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__a211o_1 _2607_ (.A1(\dataMemory[16][30] ),
    .A2(net181),
    .B1(_1755_),
    .C1(net220),
    .X(_1756_));
 sky130_fd_sc_hd__and3_1 _2608_ (.A(net293),
    .B(net255),
    .C(\dataMemory[27][30] ),
    .X(_1757_));
 sky130_fd_sc_hd__a221o_1 _2609_ (.A1(\dataMemory[24][30] ),
    .A2(net181),
    .B1(net149),
    .B2(\dataMemory[25][30] ),
    .C1(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__a211o_1 _2610_ (.A1(\dataMemory[26][30] ),
    .A2(net165),
    .B1(_1758_),
    .C1(net220),
    .X(_1759_));
 sky130_fd_sc_hd__mux4_1 _2611_ (.A0(\dataMemory[28][30] ),
    .A1(\dataMemory[29][30] ),
    .A2(\dataMemory[30][30] ),
    .A3(\dataMemory[31][30] ),
    .S0(net295),
    .S1(net257),
    .X(_1760_));
 sky130_fd_sc_hd__and3_1 _2612_ (.A(net293),
    .B(net255),
    .C(\dataMemory[7][30] ),
    .X(_1761_));
 sky130_fd_sc_hd__a221o_1 _2613_ (.A1(\dataMemory[6][30] ),
    .A2(net165),
    .B1(net149),
    .B2(\dataMemory[5][30] ),
    .C1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__a211o_1 _2614_ (.A1(\dataMemory[4][30] ),
    .A2(net181),
    .B1(_1762_),
    .C1(net194),
    .X(_1763_));
 sky130_fd_sc_hd__and3_1 _2615_ (.A(net293),
    .B(net255),
    .C(\dataMemory[3][30] ),
    .X(_1764_));
 sky130_fd_sc_hd__a221o_1 _2616_ (.A1(\dataMemory[2][30] ),
    .A2(net165),
    .B1(net148),
    .B2(\dataMemory[1][30] ),
    .C1(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__a211o_1 _2617_ (.A1(\dataMemory[0][30] ),
    .A2(net181),
    .B1(_1765_),
    .C1(net220),
    .X(_1766_));
 sky130_fd_sc_hd__and3_1 _2618_ (.A(net293),
    .B(net255),
    .C(\dataMemory[11][30] ),
    .X(_1767_));
 sky130_fd_sc_hd__a221o_1 _2619_ (.A1(\dataMemory[8][30] ),
    .A2(net180),
    .B1(net148),
    .B2(\dataMemory[9][30] ),
    .C1(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__a211o_1 _2620_ (.A1(\dataMemory[10][30] ),
    .A2(net164),
    .B1(_1768_),
    .C1(net220),
    .X(_1769_));
 sky130_fd_sc_hd__mux4_1 _2621_ (.A0(\dataMemory[12][30] ),
    .A1(\dataMemory[13][30] ),
    .A2(\dataMemory[14][30] ),
    .A3(\dataMemory[15][30] ),
    .S0(net293),
    .S1(net255),
    .X(_1770_));
 sky130_fd_sc_hd__o21a_1 _2622_ (.A1(net194),
    .A2(_1770_),
    .B1(net210),
    .X(_1771_));
 sky130_fd_sc_hd__a32o_1 _2623_ (.A1(net185),
    .A2(_1763_),
    .A3(_1766_),
    .B1(_1769_),
    .B2(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__o21a_1 _2624_ (.A1(net194),
    .A2(_1760_),
    .B1(net210),
    .X(_1773_));
 sky130_fd_sc_hd__a32o_1 _2625_ (.A1(net185),
    .A2(_1753_),
    .A3(_1756_),
    .B1(_1759_),
    .B2(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__mux2_1 _2626_ (.A0(_1772_),
    .A1(_1774_),
    .S(net204),
    .X(net63));
 sky130_fd_sc_hd__and3_1 _2627_ (.A(net294),
    .B(net256),
    .C(\dataMemory[23][31] ),
    .X(_1775_));
 sky130_fd_sc_hd__a221o_1 _2628_ (.A1(\dataMemory[22][31] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[21][31] ),
    .C1(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__a211o_1 _2629_ (.A1(\dataMemory[20][31] ),
    .A2(net180),
    .B1(_1776_),
    .C1(net194),
    .X(_1777_));
 sky130_fd_sc_hd__and3_1 _2630_ (.A(net295),
    .B(net257),
    .C(\dataMemory[19][31] ),
    .X(_1778_));
 sky130_fd_sc_hd__a221o_1 _2631_ (.A1(\dataMemory[18][31] ),
    .A2(net165),
    .B1(net149),
    .B2(\dataMemory[17][31] ),
    .C1(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__a211o_1 _2632_ (.A1(\dataMemory[16][31] ),
    .A2(net180),
    .B1(_1779_),
    .C1(net220),
    .X(_1780_));
 sky130_fd_sc_hd__and3_1 _2633_ (.A(net294),
    .B(net256),
    .C(\dataMemory[27][31] ),
    .X(_1781_));
 sky130_fd_sc_hd__a221o_1 _2634_ (.A1(\dataMemory[24][31] ),
    .A2(net181),
    .B1(net149),
    .B2(\dataMemory[25][31] ),
    .C1(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__a211o_1 _2635_ (.A1(\dataMemory[26][31] ),
    .A2(net164),
    .B1(_1782_),
    .C1(net220),
    .X(_1783_));
 sky130_fd_sc_hd__mux4_1 _2636_ (.A0(\dataMemory[28][31] ),
    .A1(\dataMemory[29][31] ),
    .A2(\dataMemory[30][31] ),
    .A3(\dataMemory[31][31] ),
    .S0(net294),
    .S1(net256),
    .X(_1784_));
 sky130_fd_sc_hd__and3_1 _2637_ (.A(net293),
    .B(net255),
    .C(\dataMemory[7][31] ),
    .X(_1785_));
 sky130_fd_sc_hd__a221o_1 _2638_ (.A1(\dataMemory[6][31] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[5][31] ),
    .C1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__a211o_1 _2639_ (.A1(\dataMemory[4][31] ),
    .A2(net180),
    .B1(_1786_),
    .C1(net194),
    .X(_1787_));
 sky130_fd_sc_hd__and3_1 _2640_ (.A(net293),
    .B(net255),
    .C(\dataMemory[3][31] ),
    .X(_1788_));
 sky130_fd_sc_hd__a221o_1 _2641_ (.A1(\dataMemory[2][31] ),
    .A2(net164),
    .B1(net148),
    .B2(\dataMemory[1][31] ),
    .C1(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__a211o_1 _2642_ (.A1(\dataMemory[0][31] ),
    .A2(net180),
    .B1(_1789_),
    .C1(net221),
    .X(_1790_));
 sky130_fd_sc_hd__and3_1 _2643_ (.A(net293),
    .B(net255),
    .C(\dataMemory[11][31] ),
    .X(_1791_));
 sky130_fd_sc_hd__a221o_1 _2644_ (.A1(\dataMemory[8][31] ),
    .A2(net180),
    .B1(net148),
    .B2(\dataMemory[9][31] ),
    .C1(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__a211o_1 _2645_ (.A1(\dataMemory[10][31] ),
    .A2(net164),
    .B1(_1792_),
    .C1(net221),
    .X(_1793_));
 sky130_fd_sc_hd__mux4_1 _2646_ (.A0(\dataMemory[12][31] ),
    .A1(\dataMemory[13][31] ),
    .A2(\dataMemory[14][31] ),
    .A3(\dataMemory[15][31] ),
    .S0(net294),
    .S1(net256),
    .X(_1794_));
 sky130_fd_sc_hd__o21a_1 _2647_ (.A1(net194),
    .A2(_1794_),
    .B1(net210),
    .X(_1795_));
 sky130_fd_sc_hd__a32o_1 _2648_ (.A1(net185),
    .A2(_1787_),
    .A3(_1790_),
    .B1(_1793_),
    .B2(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__o21a_1 _2649_ (.A1(net194),
    .A2(_1784_),
    .B1(net210),
    .X(_1797_));
 sky130_fd_sc_hd__a32o_1 _2650_ (.A1(net185),
    .A2(_1777_),
    .A3(_1780_),
    .B1(_1783_),
    .B2(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__mux2_2 _2651_ (.A0(_1796_),
    .A1(_1798_),
    .S(net205),
    .X(net64));
 sky130_fd_sc_hd__and3b_2 _2652_ (.A_N(net205),
    .B(net208),
    .C(net218),
    .X(_1799_));
 sky130_fd_sc_hd__and2_1 _2653_ (.A(net39),
    .B(net162),
    .X(_1800_));
 sky130_fd_sc_hd__nand2_2 _2654_ (.A(net39),
    .B(net162),
    .Y(_1801_));
 sky130_fd_sc_hd__nand2_2 _2655_ (.A(_1799_),
    .B(_1800_),
    .Y(_1802_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(net305),
    .A1(\dataMemory[14][17] ),
    .S(_1802_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(net302),
    .A1(\dataMemory[14][18] ),
    .S(net125),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(net301),
    .A1(\dataMemory[14][19] ),
    .S(net124),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(net296),
    .A1(\dataMemory[14][20] ),
    .S(net124),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(net276),
    .A1(\dataMemory[14][21] ),
    .S(net125),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(net275),
    .A1(\dataMemory[14][22] ),
    .S(net125),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(net272),
    .A1(\dataMemory[14][23] ),
    .S(net125),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(net270),
    .A1(\dataMemory[14][24] ),
    .S(net125),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _2664_ (.A0(net268),
    .A1(\dataMemory[14][25] ),
    .S(net125),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(net267),
    .A1(\dataMemory[14][26] ),
    .S(net124),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(net264),
    .A1(\dataMemory[14][27] ),
    .S(net125),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(net262),
    .A1(\dataMemory[14][28] ),
    .S(net125),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _2668_ (.A0(net261),
    .A1(\dataMemory[14][29] ),
    .S(net125),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2669_ (.A0(net239),
    .A1(\dataMemory[14][30] ),
    .S(net125),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(net236),
    .A1(\dataMemory[14][31] ),
    .S(net125),
    .X(_0014_));
 sky130_fd_sc_hd__and3_2 _2671_ (.A(net291),
    .B(net253),
    .C(net39),
    .X(_1803_));
 sky130_fd_sc_hd__nand3_4 _2672_ (.A(net291),
    .B(net253),
    .C(net39),
    .Y(_1804_));
 sky130_fd_sc_hd__nand2_2 _2673_ (.A(_1799_),
    .B(_1803_),
    .Y(_1805_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(net202),
    .A1(\dataMemory[15][0] ),
    .S(net134),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _2675_ (.A0(net299),
    .A1(\dataMemory[15][1] ),
    .S(net134),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(net258),
    .A1(\dataMemory[15][2] ),
    .S(net134),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _2677_ (.A0(net235),
    .A1(\dataMemory[15][3] ),
    .S(net134),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(net233),
    .A1(\dataMemory[15][4] ),
    .S(net134),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _2679_ (.A0(net230),
    .A1(\dataMemory[15][5] ),
    .S(net134),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(net228),
    .A1(\dataMemory[15][6] ),
    .S(net135),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _2681_ (.A0(net226),
    .A1(\dataMemory[15][7] ),
    .S(net134),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(net225),
    .A1(\dataMemory[15][8] ),
    .S(net134),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _2683_ (.A0(net222),
    .A1(\dataMemory[15][9] ),
    .S(net134),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(net200),
    .A1(\dataMemory[15][10] ),
    .S(net134),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _2685_ (.A0(net198),
    .A1(\dataMemory[15][11] ),
    .S(_1805_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(net314),
    .A1(\dataMemory[15][12] ),
    .S(net134),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _2687_ (.A0(net313),
    .A1(\dataMemory[15][13] ),
    .S(net134),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(net311),
    .A1(\dataMemory[15][14] ),
    .S(net134),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2689_ (.A0(net309),
    .A1(\dataMemory[15][15] ),
    .S(net135),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(net307),
    .A1(\dataMemory[15][16] ),
    .S(net135),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _2691_ (.A0(net305),
    .A1(\dataMemory[15][17] ),
    .S(net135),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(net302),
    .A1(\dataMemory[15][18] ),
    .S(net135),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2693_ (.A0(net301),
    .A1(\dataMemory[15][19] ),
    .S(net134),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(net296),
    .A1(\dataMemory[15][20] ),
    .S(net134),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2695_ (.A0(net276),
    .A1(\dataMemory[15][21] ),
    .S(net135),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(net275),
    .A1(\dataMemory[15][22] ),
    .S(net135),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2697_ (.A0(net273),
    .A1(\dataMemory[15][23] ),
    .S(net135),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(net270),
    .A1(\dataMemory[15][24] ),
    .S(net135),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(net268),
    .A1(\dataMemory[15][25] ),
    .S(net135),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(net267),
    .A1(\dataMemory[15][26] ),
    .S(net134),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(net264),
    .A1(\dataMemory[15][27] ),
    .S(net135),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(net262),
    .A1(\dataMemory[15][28] ),
    .S(net135),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(net261),
    .A1(\dataMemory[15][29] ),
    .S(net135),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2704_ (.A0(net239),
    .A1(\dataMemory[15][30] ),
    .S(net135),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(net236),
    .A1(\dataMemory[15][31] ),
    .S(net135),
    .X(_0046_));
 sky130_fd_sc_hd__or3b_4 _2706_ (.A(net219),
    .B(net208),
    .C_N(net205),
    .X(_1806_));
 sky130_fd_sc_hd__and2_1 _2707_ (.A(net39),
    .B(net179),
    .X(_1807_));
 sky130_fd_sc_hd__nand2_2 _2708_ (.A(net39),
    .B(net178),
    .Y(_1808_));
 sky130_fd_sc_hd__nor2_4 _2709_ (.A(_1806_),
    .B(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__mux2_1 _2710_ (.A0(\dataMemory[16][0] ),
    .A1(net201),
    .S(net122),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(\dataMemory[16][1] ),
    .A1(net298),
    .S(net122),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2712_ (.A0(\dataMemory[16][2] ),
    .A1(net259),
    .S(net122),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(\dataMemory[16][3] ),
    .A1(net234),
    .S(net122),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2714_ (.A0(\dataMemory[16][4] ),
    .A1(net232),
    .S(net122),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(\dataMemory[16][5] ),
    .A1(net231),
    .S(net122),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(\dataMemory[16][6] ),
    .A1(net229),
    .S(net122),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(\dataMemory[16][7] ),
    .A1(net227),
    .S(net122),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(\dataMemory[16][8] ),
    .A1(net224),
    .S(net122),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(\dataMemory[16][9] ),
    .A1(net223),
    .S(net122),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(\dataMemory[16][10] ),
    .A1(net199),
    .S(net122),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(\dataMemory[16][11] ),
    .A1(net197),
    .S(net123),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2722_ (.A0(\dataMemory[16][12] ),
    .A1(net315),
    .S(net123),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(\dataMemory[16][13] ),
    .A1(net312),
    .S(net122),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(\dataMemory[16][14] ),
    .A1(net310),
    .S(net122),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2725_ (.A0(\dataMemory[16][15] ),
    .A1(net308),
    .S(net123),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2726_ (.A0(\dataMemory[16][16] ),
    .A1(net306),
    .S(net123),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(\dataMemory[16][17] ),
    .A1(net304),
    .S(net123),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(\dataMemory[16][18] ),
    .A1(net303),
    .S(net123),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(\dataMemory[16][19] ),
    .A1(net300),
    .S(net122),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(\dataMemory[16][20] ),
    .A1(net297),
    .S(net122),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2731_ (.A0(\dataMemory[16][21] ),
    .A1(net277),
    .S(net123),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(\dataMemory[16][22] ),
    .A1(net274),
    .S(net123),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(\dataMemory[16][23] ),
    .A1(net272),
    .S(net123),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(\dataMemory[16][24] ),
    .A1(net270),
    .S(net123),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(\dataMemory[16][25] ),
    .A1(net269),
    .S(net123),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2736_ (.A0(\dataMemory[16][26] ),
    .A1(net266),
    .S(net122),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(\dataMemory[16][27] ),
    .A1(net265),
    .S(net123),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(\dataMemory[16][28] ),
    .A1(net263),
    .S(net123),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2739_ (.A0(\dataMemory[16][29] ),
    .A1(net260),
    .S(net123),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(\dataMemory[16][30] ),
    .A1(net238),
    .S(net123),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(\dataMemory[16][31] ),
    .A1(net237),
    .S(net123),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _2742_ (.A(net39),
    .B(net146),
    .X(_1810_));
 sky130_fd_sc_hd__nand2_2 _2743_ (.A(net39),
    .B(net146),
    .Y(_1811_));
 sky130_fd_sc_hd__nor2_4 _2744_ (.A(_1806_),
    .B(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(\dataMemory[17][0] ),
    .A1(net201),
    .S(net120),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(\dataMemory[17][1] ),
    .A1(net298),
    .S(net120),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(\dataMemory[17][2] ),
    .A1(net258),
    .S(net120),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(\dataMemory[17][3] ),
    .A1(net234),
    .S(net120),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2749_ (.A0(\dataMemory[17][4] ),
    .A1(net232),
    .S(net120),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2750_ (.A0(\dataMemory[17][5] ),
    .A1(net231),
    .S(net120),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(\dataMemory[17][6] ),
    .A1(net229),
    .S(net120),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(\dataMemory[17][7] ),
    .A1(net227),
    .S(net120),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(\dataMemory[17][8] ),
    .A1(net224),
    .S(net120),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(\dataMemory[17][9] ),
    .A1(net223),
    .S(net120),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2755_ (.A0(\dataMemory[17][10] ),
    .A1(net199),
    .S(net120),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2756_ (.A0(\dataMemory[17][11] ),
    .A1(net197),
    .S(net121),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(\dataMemory[17][12] ),
    .A1(net315),
    .S(net121),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2758_ (.A0(\dataMemory[17][13] ),
    .A1(net312),
    .S(net120),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(\dataMemory[17][14] ),
    .A1(net310),
    .S(net120),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2760_ (.A0(\dataMemory[17][15] ),
    .A1(net308),
    .S(net121),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(\dataMemory[17][16] ),
    .A1(net306),
    .S(net121),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2762_ (.A0(\dataMemory[17][17] ),
    .A1(net304),
    .S(net121),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(\dataMemory[17][18] ),
    .A1(net303),
    .S(net121),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2764_ (.A0(\dataMemory[17][19] ),
    .A1(net300),
    .S(net120),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(\dataMemory[17][20] ),
    .A1(net297),
    .S(net120),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(\dataMemory[17][21] ),
    .A1(net277),
    .S(net121),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(\dataMemory[17][22] ),
    .A1(net274),
    .S(net121),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(\dataMemory[17][23] ),
    .A1(net272),
    .S(net121),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(\dataMemory[17][24] ),
    .A1(net270),
    .S(net121),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(\dataMemory[17][25] ),
    .A1(net269),
    .S(net121),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(\dataMemory[17][26] ),
    .A1(net266),
    .S(net120),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(\dataMemory[17][27] ),
    .A1(net265),
    .S(net121),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2773_ (.A0(\dataMemory[17][28] ),
    .A1(net263),
    .S(net121),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(\dataMemory[17][29] ),
    .A1(net260),
    .S(net121),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2775_ (.A0(\dataMemory[17][30] ),
    .A1(net238),
    .S(net121),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2776_ (.A0(\dataMemory[17][31] ),
    .A1(net237),
    .S(net121),
    .X(_0110_));
 sky130_fd_sc_hd__nor2_4 _2777_ (.A(_1801_),
    .B(_1806_),
    .Y(_1813_));
 sky130_fd_sc_hd__mux2_1 _2778_ (.A0(\dataMemory[18][0] ),
    .A1(net201),
    .S(net118),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\dataMemory[18][1] ),
    .A1(net298),
    .S(net118),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2780_ (.A0(\dataMemory[18][2] ),
    .A1(net258),
    .S(net118),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\dataMemory[18][3] ),
    .A1(net234),
    .S(net118),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2782_ (.A0(\dataMemory[18][4] ),
    .A1(net232),
    .S(net118),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\dataMemory[18][5] ),
    .A1(net230),
    .S(net118),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(\dataMemory[18][6] ),
    .A1(net229),
    .S(net118),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(\dataMemory[18][7] ),
    .A1(net227),
    .S(net118),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _2786_ (.A0(\dataMemory[18][8] ),
    .A1(net224),
    .S(net118),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(\dataMemory[18][9] ),
    .A1(net222),
    .S(net118),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2788_ (.A0(\dataMemory[18][10] ),
    .A1(net199),
    .S(net118),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(\dataMemory[18][11] ),
    .A1(net197),
    .S(net119),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(\dataMemory[18][12] ),
    .A1(net315),
    .S(net119),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(\dataMemory[18][13] ),
    .A1(net312),
    .S(net118),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\dataMemory[18][14] ),
    .A1(net310),
    .S(net118),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2793_ (.A0(\dataMemory[18][15] ),
    .A1(net308),
    .S(net119),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(\dataMemory[18][16] ),
    .A1(net306),
    .S(net119),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _2795_ (.A0(\dataMemory[18][17] ),
    .A1(net304),
    .S(net119),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\dataMemory[18][18] ),
    .A1(net303),
    .S(net119),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(\dataMemory[18][19] ),
    .A1(net300),
    .S(net118),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(\dataMemory[18][20] ),
    .A1(net297),
    .S(net118),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2799_ (.A0(\dataMemory[18][21] ),
    .A1(net277),
    .S(net119),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\dataMemory[18][22] ),
    .A1(net274),
    .S(net119),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2801_ (.A0(\dataMemory[18][23] ),
    .A1(net272),
    .S(net119),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(\dataMemory[18][24] ),
    .A1(net270),
    .S(net119),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(\dataMemory[18][25] ),
    .A1(net269),
    .S(net119),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2804_ (.A0(\dataMemory[18][26] ),
    .A1(net266),
    .S(net118),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\dataMemory[18][27] ),
    .A1(net265),
    .S(net119),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2806_ (.A0(\dataMemory[18][28] ),
    .A1(net263),
    .S(net119),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2807_ (.A0(\dataMemory[18][29] ),
    .A1(net260),
    .S(net119),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2808_ (.A0(\dataMemory[18][30] ),
    .A1(net238),
    .S(net119),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\dataMemory[18][31] ),
    .A1(net237),
    .S(net119),
    .X(_0142_));
 sky130_fd_sc_hd__nand2_2 _2810_ (.A(net193),
    .B(_1046_),
    .Y(_1814_));
 sky130_fd_sc_hd__nor2_2 _2811_ (.A(_1811_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(\dataMemory[1][0] ),
    .A1(net202),
    .S(net116),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2813_ (.A0(\dataMemory[1][1] ),
    .A1(net299),
    .S(net116),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2814_ (.A0(\dataMemory[1][2] ),
    .A1(net258),
    .S(net116),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2815_ (.A0(\dataMemory[1][3] ),
    .A1(net235),
    .S(net116),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2816_ (.A0(\dataMemory[1][4] ),
    .A1(net232),
    .S(net116),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2817_ (.A0(\dataMemory[1][5] ),
    .A1(net230),
    .S(net116),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2818_ (.A0(\dataMemory[1][6] ),
    .A1(net228),
    .S(net116),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(\dataMemory[1][7] ),
    .A1(net226),
    .S(net116),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(\dataMemory[1][8] ),
    .A1(net225),
    .S(net116),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(\dataMemory[1][9] ),
    .A1(net222),
    .S(net116),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2822_ (.A0(\dataMemory[1][10] ),
    .A1(net199),
    .S(net117),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(\dataMemory[1][11] ),
    .A1(net198),
    .S(net117),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(\dataMemory[1][12] ),
    .A1(net314),
    .S(net116),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2825_ (.A0(\dataMemory[1][13] ),
    .A1(net313),
    .S(net116),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2826_ (.A0(\dataMemory[1][14] ),
    .A1(net310),
    .S(net116),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(\dataMemory[1][15] ),
    .A1(net308),
    .S(net117),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(\dataMemory[1][16] ),
    .A1(net307),
    .S(net117),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2829_ (.A0(\dataMemory[1][17] ),
    .A1(net305),
    .S(net117),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(\dataMemory[1][18] ),
    .A1(net302),
    .S(net116),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2831_ (.A0(\dataMemory[1][19] ),
    .A1(net300),
    .S(net116),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2832_ (.A0(\dataMemory[1][20] ),
    .A1(net296),
    .S(net117),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(\dataMemory[1][21] ),
    .A1(net276),
    .S(net117),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2834_ (.A0(\dataMemory[1][22] ),
    .A1(net275),
    .S(net117),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\dataMemory[1][23] ),
    .A1(net273),
    .S(net117),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(\dataMemory[1][24] ),
    .A1(net271),
    .S(net117),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(\dataMemory[1][25] ),
    .A1(net268),
    .S(_1815_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(\dataMemory[1][26] ),
    .A1(net266),
    .S(net116),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2839_ (.A0(\dataMemory[1][27] ),
    .A1(net264),
    .S(net117),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(\dataMemory[1][28] ),
    .A1(net262),
    .S(net117),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(\dataMemory[1][29] ),
    .A1(net260),
    .S(net117),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(\dataMemory[1][30] ),
    .A1(net238),
    .S(net117),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2843_ (.A0(\dataMemory[1][31] ),
    .A1(net237),
    .S(net117),
    .X(_0174_));
 sky130_fd_sc_hd__and3_2 _2844_ (.A(net218),
    .B(net185),
    .C(net205),
    .X(_1816_));
 sky130_fd_sc_hd__and2_2 _2845_ (.A(_1807_),
    .B(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(\dataMemory[20][0] ),
    .A1(net201),
    .S(net115),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(\dataMemory[20][1] ),
    .A1(net298),
    .S(net115),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(\dataMemory[20][2] ),
    .A1(net259),
    .S(net115),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(\dataMemory[20][3] ),
    .A1(net234),
    .S(net115),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2850_ (.A0(\dataMemory[20][4] ),
    .A1(net232),
    .S(net115),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\dataMemory[20][5] ),
    .A1(net231),
    .S(net115),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2852_ (.A0(\dataMemory[20][6] ),
    .A1(net229),
    .S(net115),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\dataMemory[20][7] ),
    .A1(net227),
    .S(net115),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2854_ (.A0(\dataMemory[20][8] ),
    .A1(net224),
    .S(net115),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(\dataMemory[20][9] ),
    .A1(net223),
    .S(net115),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(\dataMemory[20][10] ),
    .A1(net199),
    .S(net115),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\dataMemory[20][11] ),
    .A1(net197),
    .S(net114),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(\dataMemory[20][12] ),
    .A1(net315),
    .S(net114),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(\dataMemory[20][13] ),
    .A1(net312),
    .S(net115),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(\dataMemory[20][14] ),
    .A1(net310),
    .S(net115),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(\dataMemory[20][15] ),
    .A1(net308),
    .S(net114),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(\dataMemory[20][16] ),
    .A1(net306),
    .S(net114),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(\dataMemory[20][17] ),
    .A1(net304),
    .S(net114),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2864_ (.A0(\dataMemory[20][18] ),
    .A1(net303),
    .S(net114),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\dataMemory[20][19] ),
    .A1(net300),
    .S(net115),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2866_ (.A0(\dataMemory[20][20] ),
    .A1(net297),
    .S(net115),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(\dataMemory[20][21] ),
    .A1(net277),
    .S(net114),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2868_ (.A0(\dataMemory[20][22] ),
    .A1(net274),
    .S(net114),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(\dataMemory[20][23] ),
    .A1(net272),
    .S(net114),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2870_ (.A0(\dataMemory[20][24] ),
    .A1(net270),
    .S(net114),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(\dataMemory[20][25] ),
    .A1(net269),
    .S(_1817_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(\dataMemory[20][26] ),
    .A1(net266),
    .S(net114),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2873_ (.A0(\dataMemory[20][27] ),
    .A1(net265),
    .S(net114),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\dataMemory[20][28] ),
    .A1(net263),
    .S(net114),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2875_ (.A0(\dataMemory[20][29] ),
    .A1(net261),
    .S(net114),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\dataMemory[20][30] ),
    .A1(net239),
    .S(net114),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _2877_ (.A0(\dataMemory[20][31] ),
    .A1(net236),
    .S(net114),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_2 _2878_ (.A(_1810_),
    .B(_1816_),
    .Y(_1818_));
 sky130_fd_sc_hd__mux2_1 _2879_ (.A0(net201),
    .A1(\dataMemory[21][0] ),
    .S(net113),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(net298),
    .A1(\dataMemory[21][1] ),
    .S(net113),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(net259),
    .A1(\dataMemory[21][2] ),
    .S(net113),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2882_ (.A0(net234),
    .A1(\dataMemory[21][3] ),
    .S(net113),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2883_ (.A0(net232),
    .A1(\dataMemory[21][4] ),
    .S(net113),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _2884_ (.A0(net231),
    .A1(\dataMemory[21][5] ),
    .S(net113),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(net229),
    .A1(\dataMemory[21][6] ),
    .S(net113),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(net227),
    .A1(\dataMemory[21][7] ),
    .S(net112),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(net224),
    .A1(\dataMemory[21][8] ),
    .S(net113),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(net223),
    .A1(\dataMemory[21][9] ),
    .S(net113),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(net200),
    .A1(\dataMemory[21][10] ),
    .S(net112),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(net197),
    .A1(\dataMemory[21][11] ),
    .S(net112),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(net315),
    .A1(\dataMemory[21][12] ),
    .S(net112),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2892_ (.A0(net312),
    .A1(\dataMemory[21][13] ),
    .S(net113),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2893_ (.A0(net310),
    .A1(\dataMemory[21][14] ),
    .S(net113),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(net308),
    .A1(\dataMemory[21][15] ),
    .S(net113),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2895_ (.A0(net306),
    .A1(\dataMemory[21][16] ),
    .S(_1818_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(net304),
    .A1(\dataMemory[21][17] ),
    .S(net112),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(net303),
    .A1(\dataMemory[21][18] ),
    .S(net112),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(net300),
    .A1(\dataMemory[21][19] ),
    .S(net113),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(net297),
    .A1(\dataMemory[21][20] ),
    .S(net113),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(net277),
    .A1(\dataMemory[21][21] ),
    .S(net112),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(net274),
    .A1(\dataMemory[21][22] ),
    .S(net112),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(net272),
    .A1(\dataMemory[21][23] ),
    .S(net112),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(net270),
    .A1(\dataMemory[21][24] ),
    .S(net112),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2904_ (.A0(net268),
    .A1(\dataMemory[21][25] ),
    .S(net113),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(net266),
    .A1(\dataMemory[21][26] ),
    .S(net112),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2906_ (.A0(net265),
    .A1(\dataMemory[21][27] ),
    .S(net112),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2907_ (.A0(net263),
    .A1(\dataMemory[21][28] ),
    .S(net112),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(net261),
    .A1(\dataMemory[21][29] ),
    .S(net112),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(net239),
    .A1(\dataMemory[21][30] ),
    .S(net112),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2910_ (.A0(net236),
    .A1(\dataMemory[21][31] ),
    .S(net112),
    .X(_0238_));
 sky130_fd_sc_hd__nand2_2 _2911_ (.A(_1800_),
    .B(_1816_),
    .Y(_1819_));
 sky130_fd_sc_hd__mux2_1 _2912_ (.A0(net201),
    .A1(\dataMemory[22][0] ),
    .S(net111),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(net298),
    .A1(\dataMemory[22][1] ),
    .S(net111),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2914_ (.A0(net259),
    .A1(\dataMemory[22][2] ),
    .S(net111),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(net234),
    .A1(\dataMemory[22][3] ),
    .S(net111),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(net232),
    .A1(\dataMemory[22][4] ),
    .S(net111),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2917_ (.A0(net231),
    .A1(\dataMemory[22][5] ),
    .S(net111),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(net229),
    .A1(\dataMemory[22][6] ),
    .S(net111),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(net227),
    .A1(\dataMemory[22][7] ),
    .S(net110),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(net224),
    .A1(\dataMemory[22][8] ),
    .S(net111),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _2921_ (.A0(net223),
    .A1(\dataMemory[22][9] ),
    .S(net111),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(net200),
    .A1(\dataMemory[22][10] ),
    .S(net111),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(net197),
    .A1(\dataMemory[22][11] ),
    .S(net110),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _2924_ (.A0(net315),
    .A1(\dataMemory[22][12] ),
    .S(net110),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _2925_ (.A0(net312),
    .A1(\dataMemory[22][13] ),
    .S(net111),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2926_ (.A0(net12),
    .A1(\dataMemory[22][14] ),
    .S(net111),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(net308),
    .A1(\dataMemory[22][15] ),
    .S(net110),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(net306),
    .A1(\dataMemory[22][16] ),
    .S(net110),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(net304),
    .A1(\dataMemory[22][17] ),
    .S(net110),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2930_ (.A0(net303),
    .A1(\dataMemory[22][18] ),
    .S(net110),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(net300),
    .A1(\dataMemory[22][19] ),
    .S(net111),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(net297),
    .A1(\dataMemory[22][20] ),
    .S(net111),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(net277),
    .A1(\dataMemory[22][21] ),
    .S(net110),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(net274),
    .A1(\dataMemory[22][22] ),
    .S(net110),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _2935_ (.A0(net272),
    .A1(\dataMemory[22][23] ),
    .S(net110),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2936_ (.A0(net270),
    .A1(\dataMemory[22][24] ),
    .S(net110),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _2937_ (.A0(net268),
    .A1(\dataMemory[22][25] ),
    .S(net111),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(net266),
    .A1(\dataMemory[22][26] ),
    .S(net110),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(net265),
    .A1(\dataMemory[22][27] ),
    .S(_1819_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(net263),
    .A1(\dataMemory[22][28] ),
    .S(net110),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(net261),
    .A1(\dataMemory[22][29] ),
    .S(net110),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(net239),
    .A1(\dataMemory[22][30] ),
    .S(net110),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(net236),
    .A1(\dataMemory[22][31] ),
    .S(net110),
    .X(_0270_));
 sky130_fd_sc_hd__nand2_4 _2944_ (.A(_1803_),
    .B(_1816_),
    .Y(_1820_));
 sky130_fd_sc_hd__mux2_1 _2945_ (.A0(net201),
    .A1(\dataMemory[23][0] ),
    .S(net109),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(net298),
    .A1(\dataMemory[23][1] ),
    .S(net109),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(net259),
    .A1(\dataMemory[23][2] ),
    .S(net109),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _2948_ (.A0(net234),
    .A1(\dataMemory[23][3] ),
    .S(net109),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(net232),
    .A1(\dataMemory[23][4] ),
    .S(net109),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(net231),
    .A1(\dataMemory[23][5] ),
    .S(net109),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(net229),
    .A1(\dataMemory[23][6] ),
    .S(net109),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(net227),
    .A1(\dataMemory[23][7] ),
    .S(net108),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(net224),
    .A1(\dataMemory[23][8] ),
    .S(net109),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _2954_ (.A0(net223),
    .A1(\dataMemory[23][9] ),
    .S(net109),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(net200),
    .A1(\dataMemory[23][10] ),
    .S(net109),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(net197),
    .A1(\dataMemory[23][11] ),
    .S(net108),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(net315),
    .A1(\dataMemory[23][12] ),
    .S(net108),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(net312),
    .A1(\dataMemory[23][13] ),
    .S(net109),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(net310),
    .A1(\dataMemory[23][14] ),
    .S(net109),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(net13),
    .A1(\dataMemory[23][15] ),
    .S(net108),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(net306),
    .A1(\dataMemory[23][16] ),
    .S(net108),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(net304),
    .A1(\dataMemory[23][17] ),
    .S(net108),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _2963_ (.A0(net303),
    .A1(\dataMemory[23][18] ),
    .S(net108),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(net300),
    .A1(\dataMemory[23][19] ),
    .S(net109),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(net297),
    .A1(\dataMemory[23][20] ),
    .S(net109),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(net277),
    .A1(\dataMemory[23][21] ),
    .S(net108),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(net274),
    .A1(\dataMemory[23][22] ),
    .S(net108),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(net272),
    .A1(\dataMemory[23][23] ),
    .S(net108),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(net270),
    .A1(\dataMemory[23][24] ),
    .S(net108),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(net268),
    .A1(\dataMemory[23][25] ),
    .S(net109),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(net266),
    .A1(\dataMemory[23][26] ),
    .S(net108),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _2972_ (.A0(net265),
    .A1(\dataMemory[23][27] ),
    .S(_1820_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(net263),
    .A1(\dataMemory[23][28] ),
    .S(net108),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(net261),
    .A1(\dataMemory[23][29] ),
    .S(net108),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(net239),
    .A1(\dataMemory[23][30] ),
    .S(net108),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(net236),
    .A1(\dataMemory[23][31] ),
    .S(net108),
    .X(_0302_));
 sky130_fd_sc_hd__and3b_4 _2977_ (.A_N(_1039_),
    .B(_1807_),
    .C(net193),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(\dataMemory[24][0] ),
    .A1(net201),
    .S(net106),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(\dataMemory[24][1] ),
    .A1(net298),
    .S(net106),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(\dataMemory[24][2] ),
    .A1(net259),
    .S(net106),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2981_ (.A0(\dataMemory[24][3] ),
    .A1(net234),
    .S(net106),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(\dataMemory[24][4] ),
    .A1(net232),
    .S(net106),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(\dataMemory[24][5] ),
    .A1(net231),
    .S(net106),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(\dataMemory[24][6] ),
    .A1(net229),
    .S(net106),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(\dataMemory[24][7] ),
    .A1(net227),
    .S(net106),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(\dataMemory[24][8] ),
    .A1(net224),
    .S(net106),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(\dataMemory[24][9] ),
    .A1(net223),
    .S(net106),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(\dataMemory[24][10] ),
    .A1(net200),
    .S(net106),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(\dataMemory[24][11] ),
    .A1(net197),
    .S(net107),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(\dataMemory[24][12] ),
    .A1(net315),
    .S(net107),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(\dataMemory[24][13] ),
    .A1(net312),
    .S(net106),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(\dataMemory[24][14] ),
    .A1(net310),
    .S(net106),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(\dataMemory[24][15] ),
    .A1(net309),
    .S(net107),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(\dataMemory[24][16] ),
    .A1(net306),
    .S(net107),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(\dataMemory[24][17] ),
    .A1(net304),
    .S(net107),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(\dataMemory[24][18] ),
    .A1(net303),
    .S(net107),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(\dataMemory[24][19] ),
    .A1(net300),
    .S(net106),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(\dataMemory[24][20] ),
    .A1(net297),
    .S(net106),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(\dataMemory[24][21] ),
    .A1(net276),
    .S(net107),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(\dataMemory[24][22] ),
    .A1(net274),
    .S(net107),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(\dataMemory[24][23] ),
    .A1(net272),
    .S(net107),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(\dataMemory[24][24] ),
    .A1(net271),
    .S(net107),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(\dataMemory[24][25] ),
    .A1(net269),
    .S(net107),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3004_ (.A0(\dataMemory[24][26] ),
    .A1(net266),
    .S(net106),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(\dataMemory[24][27] ),
    .A1(net265),
    .S(net107),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _3006_ (.A0(\dataMemory[24][28] ),
    .A1(net263),
    .S(net107),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3007_ (.A0(\dataMemory[24][29] ),
    .A1(net28),
    .S(net107),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(\dataMemory[24][30] ),
    .A1(net238),
    .S(net107),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(\dataMemory[24][31] ),
    .A1(net237),
    .S(net107),
    .X(_0334_));
 sky130_fd_sc_hd__or3_4 _3010_ (.A(net218),
    .B(_1039_),
    .C(_1811_),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(net201),
    .A1(\dataMemory[25][0] ),
    .S(net104),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(net298),
    .A1(\dataMemory[25][1] ),
    .S(net104),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(net259),
    .A1(\dataMemory[25][2] ),
    .S(net104),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(net234),
    .A1(\dataMemory[25][3] ),
    .S(net104),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(net232),
    .A1(\dataMemory[25][4] ),
    .S(net104),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(net231),
    .A1(\dataMemory[25][5] ),
    .S(net104),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3017_ (.A0(net229),
    .A1(\dataMemory[25][6] ),
    .S(net104),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(net227),
    .A1(\dataMemory[25][7] ),
    .S(net104),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _3019_ (.A0(net224),
    .A1(\dataMemory[25][8] ),
    .S(net104),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(net223),
    .A1(\dataMemory[25][9] ),
    .S(net104),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3021_ (.A0(net200),
    .A1(\dataMemory[25][10] ),
    .S(net104),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(net197),
    .A1(\dataMemory[25][11] ),
    .S(net105),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(net315),
    .A1(\dataMemory[25][12] ),
    .S(net105),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(net312),
    .A1(\dataMemory[25][13] ),
    .S(net104),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _3025_ (.A0(net310),
    .A1(\dataMemory[25][14] ),
    .S(net104),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _3026_ (.A0(net309),
    .A1(\dataMemory[25][15] ),
    .S(net105),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(net306),
    .A1(\dataMemory[25][16] ),
    .S(net105),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(net304),
    .A1(\dataMemory[25][17] ),
    .S(net105),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _3029_ (.A0(net303),
    .A1(\dataMemory[25][18] ),
    .S(net105),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(net300),
    .A1(\dataMemory[25][19] ),
    .S(net104),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(net297),
    .A1(\dataMemory[25][20] ),
    .S(net104),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(net276),
    .A1(\dataMemory[25][21] ),
    .S(net105),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(net274),
    .A1(\dataMemory[25][22] ),
    .S(net105),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(net272),
    .A1(\dataMemory[25][23] ),
    .S(net105),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _3035_ (.A0(net270),
    .A1(\dataMemory[25][24] ),
    .S(net105),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(net269),
    .A1(\dataMemory[25][25] ),
    .S(net105),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _3037_ (.A0(net266),
    .A1(\dataMemory[25][26] ),
    .S(net104),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(net265),
    .A1(\dataMemory[25][27] ),
    .S(net105),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(net263),
    .A1(\dataMemory[25][28] ),
    .S(net105),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(net261),
    .A1(\dataMemory[25][29] ),
    .S(net105),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(net238),
    .A1(\dataMemory[25][30] ),
    .S(net105),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(net237),
    .A1(\dataMemory[25][31] ),
    .S(net105),
    .X(_0366_));
 sky130_fd_sc_hd__or3_4 _3043_ (.A(net218),
    .B(_1039_),
    .C(_1801_),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _3044_ (.A0(net201),
    .A1(\dataMemory[26][0] ),
    .S(net102),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(net298),
    .A1(\dataMemory[26][1] ),
    .S(net102),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(net259),
    .A1(\dataMemory[26][2] ),
    .S(net102),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(net234),
    .A1(\dataMemory[26][3] ),
    .S(net102),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(net232),
    .A1(\dataMemory[26][4] ),
    .S(net102),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(net231),
    .A1(\dataMemory[26][5] ),
    .S(net102),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(net229),
    .A1(\dataMemory[26][6] ),
    .S(net102),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(net227),
    .A1(\dataMemory[26][7] ),
    .S(net102),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(net224),
    .A1(\dataMemory[26][8] ),
    .S(net102),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(net223),
    .A1(\dataMemory[26][9] ),
    .S(net102),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(net199),
    .A1(\dataMemory[26][10] ),
    .S(net102),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(net197),
    .A1(\dataMemory[26][11] ),
    .S(net103),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(net315),
    .A1(\dataMemory[26][12] ),
    .S(net103),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _3057_ (.A0(net312),
    .A1(\dataMemory[26][13] ),
    .S(net102),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(net310),
    .A1(\dataMemory[26][14] ),
    .S(net102),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(net309),
    .A1(\dataMemory[26][15] ),
    .S(net103),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(net306),
    .A1(\dataMemory[26][16] ),
    .S(net103),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(net304),
    .A1(\dataMemory[26][17] ),
    .S(net103),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(net303),
    .A1(\dataMemory[26][18] ),
    .S(net103),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(net300),
    .A1(\dataMemory[26][19] ),
    .S(net102),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(net297),
    .A1(\dataMemory[26][20] ),
    .S(net102),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(net277),
    .A1(\dataMemory[26][21] ),
    .S(net103),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _3066_ (.A0(net274),
    .A1(\dataMemory[26][22] ),
    .S(net103),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3067_ (.A0(net272),
    .A1(\dataMemory[26][23] ),
    .S(net103),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(net270),
    .A1(\dataMemory[26][24] ),
    .S(net103),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3069_ (.A0(net269),
    .A1(\dataMemory[26][25] ),
    .S(net103),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(net266),
    .A1(\dataMemory[26][26] ),
    .S(net102),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3071_ (.A0(net265),
    .A1(\dataMemory[26][27] ),
    .S(net103),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(net263),
    .A1(\dataMemory[26][28] ),
    .S(net103),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _3073_ (.A0(net261),
    .A1(\dataMemory[26][29] ),
    .S(net103),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(net238),
    .A1(\dataMemory[26][30] ),
    .S(net103),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3075_ (.A0(net237),
    .A1(\dataMemory[26][31] ),
    .S(net103),
    .X(_0398_));
 sky130_fd_sc_hd__or3_4 _3076_ (.A(net218),
    .B(_1039_),
    .C(_1804_),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(net201),
    .A1(\dataMemory[27][0] ),
    .S(net132),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _3078_ (.A0(net298),
    .A1(\dataMemory[27][1] ),
    .S(net132),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(net259),
    .A1(\dataMemory[27][2] ),
    .S(net132),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3080_ (.A0(net234),
    .A1(\dataMemory[27][3] ),
    .S(net132),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(net232),
    .A1(\dataMemory[27][4] ),
    .S(net132),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _3082_ (.A0(net231),
    .A1(\dataMemory[27][5] ),
    .S(net132),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(net229),
    .A1(\dataMemory[27][6] ),
    .S(net132),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(net226),
    .A1(\dataMemory[27][7] ),
    .S(net132),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(net224),
    .A1(\dataMemory[27][8] ),
    .S(net132),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(net223),
    .A1(\dataMemory[27][9] ),
    .S(net132),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(net200),
    .A1(\dataMemory[27][10] ),
    .S(net132),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(net197),
    .A1(\dataMemory[27][11] ),
    .S(net133),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(net315),
    .A1(\dataMemory[27][12] ),
    .S(net133),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(net312),
    .A1(\dataMemory[27][13] ),
    .S(net132),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(net310),
    .A1(\dataMemory[27][14] ),
    .S(net132),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(net309),
    .A1(\dataMemory[27][15] ),
    .S(net133),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(net306),
    .A1(\dataMemory[27][16] ),
    .S(net133),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(net304),
    .A1(\dataMemory[27][17] ),
    .S(net133),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(net303),
    .A1(\dataMemory[27][18] ),
    .S(net133),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(net300),
    .A1(\dataMemory[27][19] ),
    .S(net132),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(net297),
    .A1(\dataMemory[27][20] ),
    .S(net132),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3098_ (.A0(net276),
    .A1(\dataMemory[27][21] ),
    .S(net133),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(net274),
    .A1(\dataMemory[27][22] ),
    .S(net133),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(net272),
    .A1(\dataMemory[27][23] ),
    .S(net133),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(net270),
    .A1(\dataMemory[27][24] ),
    .S(net133),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3102_ (.A0(net269),
    .A1(\dataMemory[27][25] ),
    .S(net133),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(net266),
    .A1(\dataMemory[27][26] ),
    .S(net132),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3104_ (.A0(net265),
    .A1(\dataMemory[27][27] ),
    .S(net133),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(net263),
    .A1(\dataMemory[27][28] ),
    .S(net133),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(net261),
    .A1(\dataMemory[27][29] ),
    .S(net133),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(net239),
    .A1(\dataMemory[27][30] ),
    .S(net133),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(net236),
    .A1(\dataMemory[27][31] ),
    .S(net133),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_2 _3109_ (.A(net193),
    .B(_1039_),
    .Y(_1825_));
 sky130_fd_sc_hd__nand2_2 _3110_ (.A(_1807_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(net201),
    .A1(\dataMemory[28][0] ),
    .S(net101),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(net298),
    .A1(\dataMemory[28][1] ),
    .S(net101),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(net259),
    .A1(\dataMemory[28][2] ),
    .S(net101),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(net234),
    .A1(\dataMemory[28][3] ),
    .S(net101),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _3115_ (.A0(net33),
    .A1(\dataMemory[28][4] ),
    .S(net101),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(net231),
    .A1(\dataMemory[28][5] ),
    .S(net101),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(net229),
    .A1(\dataMemory[28][6] ),
    .S(net101),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(net227),
    .A1(\dataMemory[28][7] ),
    .S(net101),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(net224),
    .A1(\dataMemory[28][8] ),
    .S(net101),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(net223),
    .A1(\dataMemory[28][9] ),
    .S(net101),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(net200),
    .A1(\dataMemory[28][10] ),
    .S(net101),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(net197),
    .A1(\dataMemory[28][11] ),
    .S(net100),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(net315),
    .A1(\dataMemory[28][12] ),
    .S(net100),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3124_ (.A0(net312),
    .A1(\dataMemory[28][13] ),
    .S(net101),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(net310),
    .A1(\dataMemory[28][14] ),
    .S(net101),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(net309),
    .A1(\dataMemory[28][15] ),
    .S(net100),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(net306),
    .A1(\dataMemory[28][16] ),
    .S(net100),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(net304),
    .A1(\dataMemory[28][17] ),
    .S(net100),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(net303),
    .A1(\dataMemory[28][18] ),
    .S(net100),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(net17),
    .A1(\dataMemory[28][19] ),
    .S(net101),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(net297),
    .A1(\dataMemory[28][20] ),
    .S(net101),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(net276),
    .A1(\dataMemory[28][21] ),
    .S(net100),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(net274),
    .A1(\dataMemory[28][22] ),
    .S(net100),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(net272),
    .A1(\dataMemory[28][23] ),
    .S(net100),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(net270),
    .A1(\dataMemory[28][24] ),
    .S(net100),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(net269),
    .A1(\dataMemory[28][25] ),
    .S(_1826_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(net266),
    .A1(\dataMemory[28][26] ),
    .S(net100),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(net265),
    .A1(\dataMemory[28][27] ),
    .S(net100),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(net263),
    .A1(\dataMemory[28][28] ),
    .S(net100),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(net261),
    .A1(\dataMemory[28][29] ),
    .S(net100),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(net239),
    .A1(\dataMemory[28][30] ),
    .S(net100),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(net236),
    .A1(\dataMemory[28][31] ),
    .S(net100),
    .X(_0462_));
 sky130_fd_sc_hd__nor2_2 _3143_ (.A(_1801_),
    .B(_1814_),
    .Y(_1827_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(\dataMemory[2][0] ),
    .A1(net202),
    .S(net98),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(\dataMemory[2][1] ),
    .A1(net299),
    .S(net98),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(\dataMemory[2][2] ),
    .A1(net258),
    .S(net98),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(\dataMemory[2][3] ),
    .A1(net235),
    .S(net98),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(\dataMemory[2][4] ),
    .A1(net233),
    .S(net98),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(\dataMemory[2][5] ),
    .A1(net230),
    .S(net98),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(\dataMemory[2][6] ),
    .A1(net228),
    .S(net98),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3151_ (.A0(\dataMemory[2][7] ),
    .A1(net226),
    .S(net98),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3152_ (.A0(\dataMemory[2][8] ),
    .A1(net225),
    .S(net98),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(\dataMemory[2][9] ),
    .A1(net222),
    .S(net98),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3154_ (.A0(\dataMemory[2][10] ),
    .A1(net199),
    .S(net99),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(\dataMemory[2][11] ),
    .A1(net198),
    .S(net99),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(\dataMemory[2][12] ),
    .A1(net314),
    .S(net98),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(\dataMemory[2][13] ),
    .A1(net313),
    .S(net98),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(\dataMemory[2][14] ),
    .A1(net311),
    .S(net98),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(\dataMemory[2][15] ),
    .A1(net308),
    .S(net99),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(\dataMemory[2][16] ),
    .A1(net307),
    .S(net99),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3161_ (.A0(\dataMemory[2][17] ),
    .A1(net305),
    .S(net99),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(\dataMemory[2][18] ),
    .A1(net302),
    .S(net98),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(\dataMemory[2][19] ),
    .A1(net300),
    .S(net98),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(\dataMemory[2][20] ),
    .A1(net296),
    .S(net99),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(\dataMemory[2][21] ),
    .A1(net276),
    .S(net99),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3166_ (.A0(\dataMemory[2][22] ),
    .A1(net275),
    .S(net99),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(\dataMemory[2][23] ),
    .A1(net273),
    .S(net99),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3168_ (.A0(\dataMemory[2][24] ),
    .A1(net271),
    .S(net99),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(\dataMemory[2][25] ),
    .A1(net268),
    .S(_1827_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3170_ (.A0(\dataMemory[2][26] ),
    .A1(net266),
    .S(net98),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(\dataMemory[2][27] ),
    .A1(net264),
    .S(net99),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3172_ (.A0(\dataMemory[2][28] ),
    .A1(net262),
    .S(net99),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(\dataMemory[2][29] ),
    .A1(net260),
    .S(net99),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3174_ (.A0(\dataMemory[2][30] ),
    .A1(net238),
    .S(net99),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(\dataMemory[2][31] ),
    .A1(net237),
    .S(net99),
    .X(_0494_));
 sky130_fd_sc_hd__nand2_2 _3176_ (.A(_1800_),
    .B(_1825_),
    .Y(_1828_));
 sky130_fd_sc_hd__mux2_1 _3177_ (.A0(net201),
    .A1(\dataMemory[30][0] ),
    .S(net97),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(net298),
    .A1(\dataMemory[30][1] ),
    .S(net97),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3179_ (.A0(net259),
    .A1(\dataMemory[30][2] ),
    .S(net97),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(net234),
    .A1(\dataMemory[30][3] ),
    .S(net97),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(net232),
    .A1(\dataMemory[30][4] ),
    .S(net97),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(net231),
    .A1(\dataMemory[30][5] ),
    .S(net97),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(net229),
    .A1(\dataMemory[30][6] ),
    .S(net97),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3184_ (.A0(net227),
    .A1(\dataMemory[30][7] ),
    .S(net97),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(net224),
    .A1(\dataMemory[30][8] ),
    .S(net97),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(net223),
    .A1(\dataMemory[30][9] ),
    .S(net97),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(net200),
    .A1(\dataMemory[30][10] ),
    .S(net97),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(net197),
    .A1(\dataMemory[30][11] ),
    .S(net96),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(net315),
    .A1(\dataMemory[30][12] ),
    .S(net96),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(net312),
    .A1(\dataMemory[30][13] ),
    .S(net97),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(net310),
    .A1(\dataMemory[30][14] ),
    .S(net97),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(net309),
    .A1(\dataMemory[30][15] ),
    .S(net96),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(net306),
    .A1(\dataMemory[30][16] ),
    .S(net96),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(net304),
    .A1(\dataMemory[30][17] ),
    .S(net96),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(net303),
    .A1(\dataMemory[30][18] ),
    .S(net96),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(net301),
    .A1(\dataMemory[30][19] ),
    .S(net97),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(net297),
    .A1(\dataMemory[30][20] ),
    .S(net97),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(net276),
    .A1(\dataMemory[30][21] ),
    .S(net96),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _3199_ (.A0(net274),
    .A1(\dataMemory[30][22] ),
    .S(net96),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(net272),
    .A1(\dataMemory[30][23] ),
    .S(net96),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(net270),
    .A1(\dataMemory[30][24] ),
    .S(net96),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(net269),
    .A1(\dataMemory[30][25] ),
    .S(_1828_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(net266),
    .A1(\dataMemory[30][26] ),
    .S(net96),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(net265),
    .A1(\dataMemory[30][27] ),
    .S(net96),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(net263),
    .A1(\dataMemory[30][28] ),
    .S(net96),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(net261),
    .A1(\dataMemory[30][29] ),
    .S(net96),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(net239),
    .A1(\dataMemory[30][30] ),
    .S(net96),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(net236),
    .A1(\dataMemory[30][31] ),
    .S(net96),
    .X(_0526_));
 sky130_fd_sc_hd__or3_4 _3209_ (.A(net219),
    .B(net185),
    .C(net205),
    .X(_1829_));
 sky130_fd_sc_hd__nor2_2 _3210_ (.A(_1811_),
    .B(_1829_),
    .Y(_1830_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(\dataMemory[9][0] ),
    .A1(net202),
    .S(net94),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(\dataMemory[9][1] ),
    .A1(net299),
    .S(net94),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(\dataMemory[9][2] ),
    .A1(net258),
    .S(net94),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(\dataMemory[9][3] ),
    .A1(net235),
    .S(net94),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\dataMemory[9][4] ),
    .A1(net233),
    .S(net94),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(\dataMemory[9][5] ),
    .A1(net230),
    .S(net94),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(\dataMemory[9][6] ),
    .A1(net228),
    .S(net94),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(\dataMemory[9][7] ),
    .A1(net226),
    .S(net94),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(\dataMemory[9][8] ),
    .A1(net225),
    .S(net94),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(\dataMemory[9][9] ),
    .A1(net222),
    .S(net94),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\dataMemory[9][10] ),
    .A1(net199),
    .S(net95),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(\dataMemory[9][11] ),
    .A1(net198),
    .S(net95),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\dataMemory[9][12] ),
    .A1(net314),
    .S(net94),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(\dataMemory[9][13] ),
    .A1(net313),
    .S(net94),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(\dataMemory[9][14] ),
    .A1(net311),
    .S(net94),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(\dataMemory[9][15] ),
    .A1(net308),
    .S(net95),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\dataMemory[9][16] ),
    .A1(net307),
    .S(net95),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(\dataMemory[9][17] ),
    .A1(net305),
    .S(net95),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(\dataMemory[9][18] ),
    .A1(net302),
    .S(net95),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(\dataMemory[9][19] ),
    .A1(net301),
    .S(net94),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(\dataMemory[9][20] ),
    .A1(net296),
    .S(net94),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(\dataMemory[9][21] ),
    .A1(net277),
    .S(net95),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(\dataMemory[9][22] ),
    .A1(net275),
    .S(net95),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(\dataMemory[9][23] ),
    .A1(net273),
    .S(net95),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(\dataMemory[9][24] ),
    .A1(net271),
    .S(net95),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(\dataMemory[9][25] ),
    .A1(net268),
    .S(_1830_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(\dataMemory[9][26] ),
    .A1(net267),
    .S(net94),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(\dataMemory[9][27] ),
    .A1(net264),
    .S(net95),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(\dataMemory[9][28] ),
    .A1(net262),
    .S(net95),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(\dataMemory[9][29] ),
    .A1(net260),
    .S(net95),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(\dataMemory[9][30] ),
    .A1(net238),
    .S(net95),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(\dataMemory[9][31] ),
    .A1(net236),
    .S(net95),
    .X(_0558_));
 sky130_fd_sc_hd__and3_2 _3243_ (.A(net218),
    .B(_1046_),
    .C(_1810_),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(\dataMemory[5][0] ),
    .A1(net202),
    .S(net92),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(\dataMemory[5][1] ),
    .A1(net299),
    .S(net92),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(\dataMemory[5][2] ),
    .A1(net258),
    .S(net92),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(\dataMemory[5][3] ),
    .A1(net235),
    .S(net92),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(\dataMemory[5][4] ),
    .A1(net233),
    .S(net92),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(\dataMemory[5][5] ),
    .A1(net230),
    .S(net92),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(\dataMemory[5][6] ),
    .A1(net228),
    .S(net92),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(\dataMemory[5][7] ),
    .A1(net226),
    .S(net92),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(\dataMemory[5][8] ),
    .A1(net225),
    .S(net92),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(\dataMemory[5][9] ),
    .A1(net222),
    .S(net92),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(\dataMemory[5][10] ),
    .A1(net199),
    .S(net93),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(\dataMemory[5][11] ),
    .A1(net198),
    .S(net93),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(\dataMemory[5][12] ),
    .A1(net314),
    .S(net92),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(\dataMemory[5][13] ),
    .A1(net313),
    .S(net92),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(\dataMemory[5][14] ),
    .A1(net311),
    .S(net92),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _3259_ (.A0(\dataMemory[5][15] ),
    .A1(net309),
    .S(net92),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(\dataMemory[5][16] ),
    .A1(net307),
    .S(net93),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(\dataMemory[5][17] ),
    .A1(net305),
    .S(net93),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\dataMemory[5][18] ),
    .A1(net302),
    .S(net93),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(\dataMemory[5][19] ),
    .A1(net301),
    .S(net92),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(\dataMemory[5][20] ),
    .A1(net296),
    .S(net93),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(\dataMemory[5][21] ),
    .A1(net277),
    .S(net93),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(\dataMemory[5][22] ),
    .A1(net275),
    .S(net93),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(\dataMemory[5][23] ),
    .A1(net273),
    .S(net93),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _3268_ (.A0(\dataMemory[5][24] ),
    .A1(net271),
    .S(net93),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(\dataMemory[5][25] ),
    .A1(net268),
    .S(_1831_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(\dataMemory[5][26] ),
    .A1(net267),
    .S(net92),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(\dataMemory[5][27] ),
    .A1(net264),
    .S(net93),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(\dataMemory[5][28] ),
    .A1(net262),
    .S(net93),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(\dataMemory[5][29] ),
    .A1(net260),
    .S(net93),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(\dataMemory[5][30] ),
    .A1(net238),
    .S(net93),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(\dataMemory[5][31] ),
    .A1(net237),
    .S(net93),
    .X(_0590_));
 sky130_fd_sc_hd__and3_2 _3276_ (.A(net218),
    .B(_1046_),
    .C(_1807_),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(\dataMemory[4][0] ),
    .A1(net202),
    .S(net90),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(\dataMemory[4][1] ),
    .A1(net299),
    .S(net90),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(\dataMemory[4][2] ),
    .A1(net258),
    .S(net90),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(\dataMemory[4][3] ),
    .A1(net235),
    .S(net90),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(\dataMemory[4][4] ),
    .A1(net233),
    .S(net90),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(\dataMemory[4][5] ),
    .A1(net230),
    .S(net90),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _3283_ (.A0(\dataMemory[4][6] ),
    .A1(net228),
    .S(net90),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(\dataMemory[4][7] ),
    .A1(net226),
    .S(net90),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(\dataMemory[4][8] ),
    .A1(net225),
    .S(net90),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(\dataMemory[4][9] ),
    .A1(net222),
    .S(net90),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(\dataMemory[4][10] ),
    .A1(net199),
    .S(net91),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(\dataMemory[4][11] ),
    .A1(net198),
    .S(net91),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _3289_ (.A0(\dataMemory[4][12] ),
    .A1(net314),
    .S(net90),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\dataMemory[4][13] ),
    .A1(net313),
    .S(net90),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _3291_ (.A0(\dataMemory[4][14] ),
    .A1(net311),
    .S(net90),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\dataMemory[4][15] ),
    .A1(net308),
    .S(net91),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(\dataMemory[4][16] ),
    .A1(net307),
    .S(net91),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(\dataMemory[4][17] ),
    .A1(net305),
    .S(net91),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _3295_ (.A0(\dataMemory[4][18] ),
    .A1(net302),
    .S(net91),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(\dataMemory[4][19] ),
    .A1(net301),
    .S(net90),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(\dataMemory[4][20] ),
    .A1(net296),
    .S(net90),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(\dataMemory[4][21] ),
    .A1(net277),
    .S(net91),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(\dataMemory[4][22] ),
    .A1(net275),
    .S(net91),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(\dataMemory[4][23] ),
    .A1(net273),
    .S(net91),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(\dataMemory[4][24] ),
    .A1(net271),
    .S(net91),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _3302_ (.A0(\dataMemory[4][25] ),
    .A1(net268),
    .S(_1832_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(\dataMemory[4][26] ),
    .A1(net267),
    .S(net90),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _3304_ (.A0(\dataMemory[4][27] ),
    .A1(net264),
    .S(net91),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(\dataMemory[4][28] ),
    .A1(net262),
    .S(net91),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(\dataMemory[4][29] ),
    .A1(net260),
    .S(net91),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(\dataMemory[4][30] ),
    .A1(net238),
    .S(net91),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(\dataMemory[4][31] ),
    .A1(net237),
    .S(net91),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_2 _3309_ (.A(_1804_),
    .B(_1814_),
    .Y(_1833_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(\dataMemory[3][0] ),
    .A1(net202),
    .S(net88),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(\dataMemory[3][1] ),
    .A1(net299),
    .S(net88),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(\dataMemory[3][2] ),
    .A1(net258),
    .S(net88),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(\dataMemory[3][3] ),
    .A1(net235),
    .S(net88),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(\dataMemory[3][4] ),
    .A1(net233),
    .S(net88),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\dataMemory[3][5] ),
    .A1(net230),
    .S(net88),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(\dataMemory[3][6] ),
    .A1(net228),
    .S(net88),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(\dataMemory[3][7] ),
    .A1(net226),
    .S(net88),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(\dataMemory[3][8] ),
    .A1(net225),
    .S(net88),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(\dataMemory[3][9] ),
    .A1(net222),
    .S(net88),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(\dataMemory[3][10] ),
    .A1(net199),
    .S(net89),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\dataMemory[3][11] ),
    .A1(net198),
    .S(net89),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(\dataMemory[3][12] ),
    .A1(net314),
    .S(net88),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _3323_ (.A0(\dataMemory[3][13] ),
    .A1(net313),
    .S(net88),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(\dataMemory[3][14] ),
    .A1(net311),
    .S(net88),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _3325_ (.A0(\dataMemory[3][15] ),
    .A1(net308),
    .S(net89),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _3326_ (.A0(\dataMemory[3][16] ),
    .A1(net307),
    .S(net89),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _3327_ (.A0(\dataMemory[3][17] ),
    .A1(net305),
    .S(net89),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(\dataMemory[3][18] ),
    .A1(net302),
    .S(net88),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _3329_ (.A0(\dataMemory[3][19] ),
    .A1(net300),
    .S(net88),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(\dataMemory[3][20] ),
    .A1(net296),
    .S(net89),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _3331_ (.A0(\dataMemory[3][21] ),
    .A1(net276),
    .S(net89),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(\dataMemory[3][22] ),
    .A1(net275),
    .S(net89),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _3333_ (.A0(\dataMemory[3][23] ),
    .A1(net273),
    .S(net89),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(\dataMemory[3][24] ),
    .A1(net271),
    .S(net89),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(\dataMemory[3][25] ),
    .A1(net269),
    .S(_1833_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _3336_ (.A0(\dataMemory[3][26] ),
    .A1(net266),
    .S(net88),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(\dataMemory[3][27] ),
    .A1(net264),
    .S(net89),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _3338_ (.A0(\dataMemory[3][28] ),
    .A1(net262),
    .S(net89),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(\dataMemory[3][29] ),
    .A1(net260),
    .S(net89),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(\dataMemory[3][30] ),
    .A1(net238),
    .S(net89),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _3341_ (.A0(\dataMemory[3][31] ),
    .A1(net237),
    .S(net89),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_2 _3342_ (.A(_1803_),
    .B(_1825_),
    .Y(_1834_));
 sky130_fd_sc_hd__mux2_1 _3343_ (.A0(net201),
    .A1(\dataMemory[31][0] ),
    .S(net87),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(net298),
    .A1(\dataMemory[31][1] ),
    .S(net87),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _3345_ (.A0(net259),
    .A1(\dataMemory[31][2] ),
    .S(net87),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(net234),
    .A1(\dataMemory[31][3] ),
    .S(net87),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _3347_ (.A0(net232),
    .A1(\dataMemory[31][4] ),
    .S(net87),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(net231),
    .A1(\dataMemory[31][5] ),
    .S(net87),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(net229),
    .A1(\dataMemory[31][6] ),
    .S(net87),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _3350_ (.A0(net227),
    .A1(\dataMemory[31][7] ),
    .S(net87),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(net224),
    .A1(\dataMemory[31][8] ),
    .S(net87),
    .X(_0663_));
 sky130_fd_sc_hd__mux2_1 _3352_ (.A0(net223),
    .A1(\dataMemory[31][9] ),
    .S(net87),
    .X(_0664_));
 sky130_fd_sc_hd__mux2_1 _3353_ (.A0(net200),
    .A1(\dataMemory[31][10] ),
    .S(net87),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_1 _3354_ (.A0(net197),
    .A1(\dataMemory[31][11] ),
    .S(net86),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(net315),
    .A1(\dataMemory[31][12] ),
    .S(net86),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _3356_ (.A0(net312),
    .A1(\dataMemory[31][13] ),
    .S(net87),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(net310),
    .A1(\dataMemory[31][14] ),
    .S(net87),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(net309),
    .A1(\dataMemory[31][15] ),
    .S(net86),
    .X(_0670_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(net306),
    .A1(\dataMemory[31][16] ),
    .S(net86),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_1 _3360_ (.A0(net304),
    .A1(\dataMemory[31][17] ),
    .S(net86),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(net303),
    .A1(\dataMemory[31][18] ),
    .S(net86),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _3362_ (.A0(net301),
    .A1(\dataMemory[31][19] ),
    .S(net87),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_1 _3363_ (.A0(net297),
    .A1(\dataMemory[31][20] ),
    .S(net87),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(net276),
    .A1(\dataMemory[31][21] ),
    .S(net86),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(net274),
    .A1(\dataMemory[31][22] ),
    .S(net86),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(net272),
    .A1(\dataMemory[31][23] ),
    .S(net86),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(net270),
    .A1(\dataMemory[31][24] ),
    .S(net86),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(net269),
    .A1(\dataMemory[31][25] ),
    .S(_1834_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(net25),
    .A1(\dataMemory[31][26] ),
    .S(net86),
    .X(_0681_));
 sky130_fd_sc_hd__mux2_1 _3370_ (.A0(net265),
    .A1(\dataMemory[31][27] ),
    .S(net86),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(net263),
    .A1(\dataMemory[31][28] ),
    .S(net86),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_1 _3372_ (.A0(net261),
    .A1(\dataMemory[31][29] ),
    .S(net86),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(net239),
    .A1(\dataMemory[31][30] ),
    .S(net86),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(net236),
    .A1(\dataMemory[31][31] ),
    .S(net86),
    .X(_0686_));
 sky130_fd_sc_hd__nor2_4 _3375_ (.A(_1804_),
    .B(_1806_),
    .Y(_1835_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(\dataMemory[19][0] ),
    .A1(net201),
    .S(net130),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(\dataMemory[19][1] ),
    .A1(net298),
    .S(net130),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_1 _3378_ (.A0(\dataMemory[19][2] ),
    .A1(net259),
    .S(net130),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(\dataMemory[19][3] ),
    .A1(net234),
    .S(net130),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(\dataMemory[19][4] ),
    .A1(net233),
    .S(net130),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(\dataMemory[19][5] ),
    .A1(net231),
    .S(net130),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(\dataMemory[19][6] ),
    .A1(net229),
    .S(net130),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(\dataMemory[19][7] ),
    .A1(net227),
    .S(net130),
    .X(_0694_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(\dataMemory[19][8] ),
    .A1(net224),
    .S(net130),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _3385_ (.A0(\dataMemory[19][9] ),
    .A1(net223),
    .S(net130),
    .X(_0696_));
 sky130_fd_sc_hd__mux2_1 _3386_ (.A0(\dataMemory[19][10] ),
    .A1(net8),
    .S(net130),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _3387_ (.A0(\dataMemory[19][11] ),
    .A1(net197),
    .S(net131),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _3388_ (.A0(\dataMemory[19][12] ),
    .A1(net315),
    .S(net131),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _3389_ (.A0(\dataMemory[19][13] ),
    .A1(net312),
    .S(net130),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(\dataMemory[19][14] ),
    .A1(net310),
    .S(net130),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(\dataMemory[19][15] ),
    .A1(net309),
    .S(net131),
    .X(_0702_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(\dataMemory[19][16] ),
    .A1(net306),
    .S(net131),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(\dataMemory[19][17] ),
    .A1(net304),
    .S(net131),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _3394_ (.A0(\dataMemory[19][18] ),
    .A1(net303),
    .S(net131),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(\dataMemory[19][19] ),
    .A1(net301),
    .S(net130),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(\dataMemory[19][20] ),
    .A1(net297),
    .S(net130),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _3397_ (.A0(\dataMemory[19][21] ),
    .A1(net276),
    .S(net131),
    .X(_0708_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(\dataMemory[19][22] ),
    .A1(net274),
    .S(net131),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(\dataMemory[19][23] ),
    .A1(net273),
    .S(net131),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(\dataMemory[19][24] ),
    .A1(net271),
    .S(net131),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(\dataMemory[19][25] ),
    .A1(net269),
    .S(net131),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(\dataMemory[19][26] ),
    .A1(net267),
    .S(net130),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _3403_ (.A0(\dataMemory[19][27] ),
    .A1(net265),
    .S(net131),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(\dataMemory[19][28] ),
    .A1(net263),
    .S(net131),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(\dataMemory[19][29] ),
    .A1(net261),
    .S(net131),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _3406_ (.A0(\dataMemory[19][30] ),
    .A1(net30),
    .S(net131),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _3407_ (.A0(\dataMemory[19][31] ),
    .A1(net237),
    .S(net131),
    .X(_0718_));
 sky130_fd_sc_hd__and3_2 _3408_ (.A(net218),
    .B(_1046_),
    .C(_1800_),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(\dataMemory[6][0] ),
    .A1(net202),
    .S(net84),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _3410_ (.A0(\dataMemory[6][1] ),
    .A1(net299),
    .S(net84),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(\dataMemory[6][2] ),
    .A1(net258),
    .S(net84),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(\dataMemory[6][3] ),
    .A1(net235),
    .S(net84),
    .X(_0722_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(\dataMemory[6][4] ),
    .A1(net233),
    .S(net84),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(\dataMemory[6][5] ),
    .A1(net230),
    .S(net84),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(\dataMemory[6][6] ),
    .A1(net228),
    .S(net84),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _3416_ (.A0(\dataMemory[6][7] ),
    .A1(net226),
    .S(net84),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(\dataMemory[6][8] ),
    .A1(net225),
    .S(net84),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(\dataMemory[6][9] ),
    .A1(net222),
    .S(net84),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(\dataMemory[6][10] ),
    .A1(net199),
    .S(net85),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(\dataMemory[6][11] ),
    .A1(net198),
    .S(net85),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(\dataMemory[6][12] ),
    .A1(net314),
    .S(net84),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(\dataMemory[6][13] ),
    .A1(net313),
    .S(net84),
    .X(_0732_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(\dataMemory[6][14] ),
    .A1(net311),
    .S(net84),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(\dataMemory[6][15] ),
    .A1(net308),
    .S(net84),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(\dataMemory[6][16] ),
    .A1(net307),
    .S(net85),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(\dataMemory[6][17] ),
    .A1(net305),
    .S(net85),
    .X(_0736_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(\dataMemory[6][18] ),
    .A1(net302),
    .S(net85),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(\dataMemory[6][19] ),
    .A1(net301),
    .S(net84),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(\dataMemory[6][20] ),
    .A1(net296),
    .S(net85),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(\dataMemory[6][21] ),
    .A1(net277),
    .S(net85),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(\dataMemory[6][22] ),
    .A1(net275),
    .S(net85),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(\dataMemory[6][23] ),
    .A1(net273),
    .S(net85),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(\dataMemory[6][24] ),
    .A1(net271),
    .S(net85),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(\dataMemory[6][25] ),
    .A1(net269),
    .S(_1836_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(\dataMemory[6][26] ),
    .A1(net267),
    .S(net84),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(\dataMemory[6][27] ),
    .A1(net264),
    .S(net85),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _3437_ (.A0(\dataMemory[6][28] ),
    .A1(net262),
    .S(net85),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(\dataMemory[6][29] ),
    .A1(net260),
    .S(net85),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(\dataMemory[6][30] ),
    .A1(net238),
    .S(net85),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(\dataMemory[6][31] ),
    .A1(net237),
    .S(net85),
    .X(_0750_));
 sky130_fd_sc_hd__nand2_2 _3441_ (.A(_1810_),
    .B(_1825_),
    .Y(_1837_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(net201),
    .A1(\dataMemory[29][0] ),
    .S(net83),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(net298),
    .A1(\dataMemory[29][1] ),
    .S(net83),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(net259),
    .A1(\dataMemory[29][2] ),
    .S(net83),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(net234),
    .A1(\dataMemory[29][3] ),
    .S(net83),
    .X(_0754_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(net232),
    .A1(\dataMemory[29][4] ),
    .S(net83),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(net231),
    .A1(\dataMemory[29][5] ),
    .S(net83),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(net229),
    .A1(\dataMemory[29][6] ),
    .S(net83),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(net36),
    .A1(\dataMemory[29][7] ),
    .S(net83),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(net224),
    .A1(\dataMemory[29][8] ),
    .S(net83),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(net223),
    .A1(\dataMemory[29][9] ),
    .S(net83),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(net200),
    .A1(\dataMemory[29][10] ),
    .S(net83),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(net197),
    .A1(\dataMemory[29][11] ),
    .S(net82),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(net315),
    .A1(\dataMemory[29][12] ),
    .S(net82),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(net312),
    .A1(\dataMemory[29][13] ),
    .S(net83),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _3456_ (.A0(net310),
    .A1(\dataMemory[29][14] ),
    .S(net83),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(net309),
    .A1(\dataMemory[29][15] ),
    .S(net82),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(net306),
    .A1(\dataMemory[29][16] ),
    .S(net82),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _3459_ (.A0(net304),
    .A1(\dataMemory[29][17] ),
    .S(net82),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(net303),
    .A1(\dataMemory[29][18] ),
    .S(net82),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(net301),
    .A1(\dataMemory[29][19] ),
    .S(net83),
    .X(_0770_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(net297),
    .A1(\dataMemory[29][20] ),
    .S(net83),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(net276),
    .A1(\dataMemory[29][21] ),
    .S(net82),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(net274),
    .A1(\dataMemory[29][22] ),
    .S(net82),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(net272),
    .A1(\dataMemory[29][23] ),
    .S(net82),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(net270),
    .A1(\dataMemory[29][24] ),
    .S(net82),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(net24),
    .A1(\dataMemory[29][25] ),
    .S(_1837_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(net267),
    .A1(\dataMemory[29][26] ),
    .S(net82),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(net265),
    .A1(\dataMemory[29][27] ),
    .S(net82),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(net263),
    .A1(\dataMemory[29][28] ),
    .S(net82),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(net261),
    .A1(\dataMemory[29][29] ),
    .S(net82),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _3472_ (.A0(net239),
    .A1(\dataMemory[29][30] ),
    .S(net82),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(net236),
    .A1(\dataMemory[29][31] ),
    .S(net82),
    .X(_0782_));
 sky130_fd_sc_hd__and3_2 _3474_ (.A(net218),
    .B(_1046_),
    .C(_1803_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _3475_ (.A0(\dataMemory[7][0] ),
    .A1(net202),
    .S(net128),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(\dataMemory[7][1] ),
    .A1(net299),
    .S(net128),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(\dataMemory[7][2] ),
    .A1(net258),
    .S(net128),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(\dataMemory[7][3] ),
    .A1(net235),
    .S(net128),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _3479_ (.A0(\dataMemory[7][4] ),
    .A1(net233),
    .S(net128),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\dataMemory[7][5] ),
    .A1(net230),
    .S(net128),
    .X(_0788_));
 sky130_fd_sc_hd__mux2_1 _3481_ (.A0(\dataMemory[7][6] ),
    .A1(net228),
    .S(net128),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(\dataMemory[7][7] ),
    .A1(net226),
    .S(net128),
    .X(_0790_));
 sky130_fd_sc_hd__mux2_1 _3483_ (.A0(\dataMemory[7][8] ),
    .A1(net225),
    .S(net128),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(\dataMemory[7][9] ),
    .A1(net222),
    .S(net128),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(\dataMemory[7][10] ),
    .A1(net199),
    .S(net129),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(\dataMemory[7][11] ),
    .A1(net198),
    .S(net129),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(\dataMemory[7][12] ),
    .A1(net314),
    .S(net128),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(\dataMemory[7][13] ),
    .A1(net313),
    .S(net128),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(\dataMemory[7][14] ),
    .A1(net311),
    .S(net128),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(\dataMemory[7][15] ),
    .A1(net309),
    .S(net128),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _3491_ (.A0(\dataMemory[7][16] ),
    .A1(net307),
    .S(net129),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(\dataMemory[7][17] ),
    .A1(net305),
    .S(net129),
    .X(_0800_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(\dataMemory[7][18] ),
    .A1(net302),
    .S(net129),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(\dataMemory[7][19] ),
    .A1(net301),
    .S(net128),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _3495_ (.A0(\dataMemory[7][20] ),
    .A1(net296),
    .S(net129),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(\dataMemory[7][21] ),
    .A1(net277),
    .S(net129),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _3497_ (.A0(\dataMemory[7][22] ),
    .A1(net275),
    .S(net129),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(\dataMemory[7][23] ),
    .A1(net273),
    .S(net129),
    .X(_0806_));
 sky130_fd_sc_hd__mux2_1 _3499_ (.A0(\dataMemory[7][24] ),
    .A1(net271),
    .S(net129),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\dataMemory[7][25] ),
    .A1(net268),
    .S(_1838_),
    .X(_0808_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(\dataMemory[7][26] ),
    .A1(net267),
    .S(net128),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(\dataMemory[7][27] ),
    .A1(net264),
    .S(net129),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _3503_ (.A0(\dataMemory[7][28] ),
    .A1(net262),
    .S(net129),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(\dataMemory[7][29] ),
    .A1(net260),
    .S(net129),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(\dataMemory[7][30] ),
    .A1(net238),
    .S(net129),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(\dataMemory[7][31] ),
    .A1(net237),
    .S(net129),
    .X(_0814_));
 sky130_fd_sc_hd__nor2_2 _3507_ (.A(_1808_),
    .B(_1829_),
    .Y(_1839_));
 sky130_fd_sc_hd__mux2_1 _3508_ (.A0(\dataMemory[8][0] ),
    .A1(net202),
    .S(net80),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(\dataMemory[8][1] ),
    .A1(net299),
    .S(net80),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(\dataMemory[8][2] ),
    .A1(net258),
    .S(net80),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(\dataMemory[8][3] ),
    .A1(net235),
    .S(net80),
    .X(_0818_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(\dataMemory[8][4] ),
    .A1(net233),
    .S(net80),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(\dataMemory[8][5] ),
    .A1(net230),
    .S(net80),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(\dataMemory[8][6] ),
    .A1(net228),
    .S(net80),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(\dataMemory[8][7] ),
    .A1(net226),
    .S(net80),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(\dataMemory[8][8] ),
    .A1(net225),
    .S(net80),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _3517_ (.A0(\dataMemory[8][9] ),
    .A1(net222),
    .S(net80),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(\dataMemory[8][10] ),
    .A1(net199),
    .S(net81),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(\dataMemory[8][11] ),
    .A1(net198),
    .S(net81),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(\dataMemory[8][12] ),
    .A1(net314),
    .S(net80),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(\dataMemory[8][13] ),
    .A1(net313),
    .S(net80),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(\dataMemory[8][14] ),
    .A1(net311),
    .S(net80),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(\dataMemory[8][15] ),
    .A1(net308),
    .S(net81),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _3524_ (.A0(\dataMemory[8][16] ),
    .A1(net307),
    .S(net81),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(\dataMemory[8][17] ),
    .A1(net305),
    .S(net81),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(\dataMemory[8][18] ),
    .A1(net302),
    .S(net81),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _3527_ (.A0(\dataMemory[8][19] ),
    .A1(net301),
    .S(net80),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(\dataMemory[8][20] ),
    .A1(net296),
    .S(net80),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(\dataMemory[8][21] ),
    .A1(net277),
    .S(net81),
    .X(_0836_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(\dataMemory[8][22] ),
    .A1(net275),
    .S(net81),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(\dataMemory[8][23] ),
    .A1(net273),
    .S(net81),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(\dataMemory[8][24] ),
    .A1(net271),
    .S(net81),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(\dataMemory[8][25] ),
    .A1(net268),
    .S(_1839_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(\dataMemory[8][26] ),
    .A1(net267),
    .S(net80),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _3535_ (.A0(\dataMemory[8][27] ),
    .A1(net264),
    .S(net81),
    .X(_0842_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(\dataMemory[8][28] ),
    .A1(net262),
    .S(net81),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(\dataMemory[8][29] ),
    .A1(net260),
    .S(net81),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(\dataMemory[8][30] ),
    .A1(net238),
    .S(net81),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(\dataMemory[8][31] ),
    .A1(net236),
    .S(net81),
    .X(_0846_));
 sky130_fd_sc_hd__nor2_2 _3540_ (.A(_1808_),
    .B(_1814_),
    .Y(_1840_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(\dataMemory[0][0] ),
    .A1(net202),
    .S(net78),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(\dataMemory[0][1] ),
    .A1(net299),
    .S(net78),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(\dataMemory[0][2] ),
    .A1(net258),
    .S(net78),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(\dataMemory[0][3] ),
    .A1(net235),
    .S(net78),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(\dataMemory[0][4] ),
    .A1(net233),
    .S(net78),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(\dataMemory[0][5] ),
    .A1(net230),
    .S(net78),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _3547_ (.A0(\dataMemory[0][6] ),
    .A1(net228),
    .S(net78),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(\dataMemory[0][7] ),
    .A1(net226),
    .S(net78),
    .X(_0854_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(\dataMemory[0][8] ),
    .A1(net225),
    .S(net78),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\dataMemory[0][9] ),
    .A1(net222),
    .S(net78),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(\dataMemory[0][10] ),
    .A1(net199),
    .S(net79),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(\dataMemory[0][11] ),
    .A1(net198),
    .S(net79),
    .X(_0858_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(\dataMemory[0][12] ),
    .A1(net314),
    .S(net78),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(\dataMemory[0][13] ),
    .A1(net313),
    .S(net78),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(\dataMemory[0][14] ),
    .A1(net311),
    .S(net78),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(\dataMemory[0][15] ),
    .A1(net308),
    .S(net79),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\dataMemory[0][16] ),
    .A1(net307),
    .S(net79),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(\dataMemory[0][17] ),
    .A1(net305),
    .S(net79),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\dataMemory[0][18] ),
    .A1(net302),
    .S(net79),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(\dataMemory[0][19] ),
    .A1(net300),
    .S(net78),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(\dataMemory[0][20] ),
    .A1(net296),
    .S(net78),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(\dataMemory[0][21] ),
    .A1(net276),
    .S(net79),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(\dataMemory[0][22] ),
    .A1(net275),
    .S(net79),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(\dataMemory[0][23] ),
    .A1(net273),
    .S(net79),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(\dataMemory[0][24] ),
    .A1(net271),
    .S(net79),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(\dataMemory[0][25] ),
    .A1(net269),
    .S(_1840_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(\dataMemory[0][26] ),
    .A1(net267),
    .S(net78),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(\dataMemory[0][27] ),
    .A1(net264),
    .S(net79),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(\dataMemory[0][28] ),
    .A1(net262),
    .S(net79),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\dataMemory[0][29] ),
    .A1(net260),
    .S(net79),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _3571_ (.A0(\dataMemory[0][30] ),
    .A1(net239),
    .S(net79),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(\dataMemory[0][31] ),
    .A1(net237),
    .S(net79),
    .X(_0878_));
 sky130_fd_sc_hd__nor2_2 _3573_ (.A(_1801_),
    .B(_1829_),
    .Y(_1841_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\dataMemory[10][0] ),
    .A1(net202),
    .S(net76),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(\dataMemory[10][1] ),
    .A1(net299),
    .S(net76),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(\dataMemory[10][2] ),
    .A1(net29),
    .S(net76),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(\dataMemory[10][3] ),
    .A1(net235),
    .S(net76),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\dataMemory[10][4] ),
    .A1(net233),
    .S(net76),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(\dataMemory[10][5] ),
    .A1(net230),
    .S(net76),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(\dataMemory[10][6] ),
    .A1(net228),
    .S(net77),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(\dataMemory[10][7] ),
    .A1(net226),
    .S(net76),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(\dataMemory[10][8] ),
    .A1(net225),
    .S(net76),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _3583_ (.A0(\dataMemory[10][9] ),
    .A1(net38),
    .S(net76),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(\dataMemory[10][10] ),
    .A1(net199),
    .S(net76),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(\dataMemory[10][11] ),
    .A1(net198),
    .S(_1841_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(\dataMemory[10][12] ),
    .A1(net314),
    .S(net76),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _3587_ (.A0(\dataMemory[10][13] ),
    .A1(net313),
    .S(net76),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(\dataMemory[10][14] ),
    .A1(net311),
    .S(net76),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _3589_ (.A0(\dataMemory[10][15] ),
    .A1(net308),
    .S(net77),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(\dataMemory[10][16] ),
    .A1(net307),
    .S(net77),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _3591_ (.A0(\dataMemory[10][17] ),
    .A1(net305),
    .S(net77),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(\dataMemory[10][18] ),
    .A1(net302),
    .S(net77),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(\dataMemory[10][19] ),
    .A1(net301),
    .S(net76),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(\dataMemory[10][20] ),
    .A1(net296),
    .S(net76),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(\dataMemory[10][21] ),
    .A1(net277),
    .S(net77),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _3596_ (.A0(\dataMemory[10][22] ),
    .A1(net275),
    .S(net77),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(\dataMemory[10][23] ),
    .A1(net273),
    .S(net77),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _3598_ (.A0(\dataMemory[10][24] ),
    .A1(net271),
    .S(net77),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(\dataMemory[10][25] ),
    .A1(net268),
    .S(net77),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _3600_ (.A0(\dataMemory[10][26] ),
    .A1(net267),
    .S(net76),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(\dataMemory[10][27] ),
    .A1(net264),
    .S(net77),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _3602_ (.A0(\dataMemory[10][28] ),
    .A1(net262),
    .S(net77),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _3603_ (.A0(\dataMemory[10][29] ),
    .A1(net260),
    .S(net77),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _3604_ (.A0(\dataMemory[10][30] ),
    .A1(net238),
    .S(net77),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(\dataMemory[10][31] ),
    .A1(net237),
    .S(net77),
    .X(_0910_));
 sky130_fd_sc_hd__nor2_2 _3606_ (.A(_1804_),
    .B(_1829_),
    .Y(_1842_));
 sky130_fd_sc_hd__mux2_1 _3607_ (.A0(\dataMemory[11][0] ),
    .A1(net202),
    .S(net74),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(\dataMemory[11][1] ),
    .A1(net299),
    .S(net74),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _3609_ (.A0(\dataMemory[11][2] ),
    .A1(net258),
    .S(net74),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _3610_ (.A0(\dataMemory[11][3] ),
    .A1(net235),
    .S(net74),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(\dataMemory[11][4] ),
    .A1(net232),
    .S(net74),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(\dataMemory[11][5] ),
    .A1(net230),
    .S(net74),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _3613_ (.A0(\dataMemory[11][6] ),
    .A1(net228),
    .S(net74),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _3614_ (.A0(\dataMemory[11][7] ),
    .A1(net226),
    .S(net74),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _3615_ (.A0(\dataMemory[11][8] ),
    .A1(net225),
    .S(net74),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_1 _3616_ (.A0(\dataMemory[11][9] ),
    .A1(net222),
    .S(net74),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(\dataMemory[11][10] ),
    .A1(net200),
    .S(net75),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _3618_ (.A0(\dataMemory[11][11] ),
    .A1(net198),
    .S(net75),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _3619_ (.A0(\dataMemory[11][12] ),
    .A1(net314),
    .S(net74),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _3620_ (.A0(\dataMemory[11][13] ),
    .A1(net313),
    .S(net74),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(\dataMemory[11][14] ),
    .A1(net311),
    .S(net74),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _3622_ (.A0(\dataMemory[11][15] ),
    .A1(net308),
    .S(net75),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _3623_ (.A0(\dataMemory[11][16] ),
    .A1(net307),
    .S(net75),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3624_ (.A0(\dataMemory[11][17] ),
    .A1(net305),
    .S(net75),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _3625_ (.A0(\dataMemory[11][18] ),
    .A1(net302),
    .S(net75),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_1 _3626_ (.A0(\dataMemory[11][19] ),
    .A1(net301),
    .S(net74),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _3627_ (.A0(\dataMemory[11][20] ),
    .A1(net296),
    .S(net74),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _3628_ (.A0(\dataMemory[11][21] ),
    .A1(net277),
    .S(net75),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(\dataMemory[11][22] ),
    .A1(net275),
    .S(net75),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _3630_ (.A0(\dataMemory[11][23] ),
    .A1(net273),
    .S(net75),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _3631_ (.A0(\dataMemory[11][24] ),
    .A1(net271),
    .S(net75),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _3632_ (.A0(\dataMemory[11][25] ),
    .A1(net268),
    .S(_1842_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(\dataMemory[11][26] ),
    .A1(net267),
    .S(net74),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _3634_ (.A0(\dataMemory[11][27] ),
    .A1(net264),
    .S(net75),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _3635_ (.A0(\dataMemory[11][28] ),
    .A1(net262),
    .S(net75),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(\dataMemory[11][29] ),
    .A1(net260),
    .S(net75),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(\dataMemory[11][30] ),
    .A1(net239),
    .S(net75),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _3638_ (.A0(\dataMemory[11][31] ),
    .A1(net236),
    .S(net75),
    .X(_0942_));
 sky130_fd_sc_hd__and3_2 _3639_ (.A(net39),
    .B(net179),
    .C(_1799_),
    .X(_1843_));
 sky130_fd_sc_hd__mux2_1 _3640_ (.A0(\dataMemory[12][0] ),
    .A1(net202),
    .S(net126),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _3641_ (.A0(\dataMemory[12][1] ),
    .A1(net299),
    .S(net126),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _3642_ (.A0(\dataMemory[12][2] ),
    .A1(net259),
    .S(net126),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _3643_ (.A0(\dataMemory[12][3] ),
    .A1(net235),
    .S(net126),
    .X(_0946_));
 sky130_fd_sc_hd__mux2_1 _3644_ (.A0(\dataMemory[12][4] ),
    .A1(net233),
    .S(net126),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(\dataMemory[12][5] ),
    .A1(net34),
    .S(net126),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _3646_ (.A0(\dataMemory[12][6] ),
    .A1(net228),
    .S(net126),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _3647_ (.A0(\dataMemory[12][7] ),
    .A1(net226),
    .S(net127),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _3648_ (.A0(\dataMemory[12][8] ),
    .A1(net225),
    .S(net126),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(\dataMemory[12][9] ),
    .A1(net222),
    .S(net126),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(\dataMemory[12][10] ),
    .A1(net200),
    .S(net126),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _3651_ (.A0(\dataMemory[12][11] ),
    .A1(net198),
    .S(_1843_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(\dataMemory[12][12] ),
    .A1(net314),
    .S(net126),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(\dataMemory[12][13] ),
    .A1(net313),
    .S(net126),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3654_ (.A0(\dataMemory[12][14] ),
    .A1(net311),
    .S(net126),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3655_ (.A0(\dataMemory[12][15] ),
    .A1(net309),
    .S(net127),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3656_ (.A0(\dataMemory[12][16] ),
    .A1(net307),
    .S(net127),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(\dataMemory[12][17] ),
    .A1(net305),
    .S(net127),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(\dataMemory[12][18] ),
    .A1(net302),
    .S(net127),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(\dataMemory[12][19] ),
    .A1(net301),
    .S(net126),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\dataMemory[12][20] ),
    .A1(net296),
    .S(net126),
    .X(_0963_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(\dataMemory[12][21] ),
    .A1(net276),
    .S(net127),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(\dataMemory[12][22] ),
    .A1(net275),
    .S(net127),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(\dataMemory[12][23] ),
    .A1(net273),
    .S(net127),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(\dataMemory[12][24] ),
    .A1(net23),
    .S(net127),
    .X(_0967_));
 sky130_fd_sc_hd__mux2_1 _3665_ (.A0(\dataMemory[12][25] ),
    .A1(net268),
    .S(net127),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(\dataMemory[12][26] ),
    .A1(net267),
    .S(net126),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(\dataMemory[12][27] ),
    .A1(net264),
    .S(net127),
    .X(_0970_));
 sky130_fd_sc_hd__mux2_1 _3668_ (.A0(\dataMemory[12][28] ),
    .A1(net262),
    .S(net127),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(\dataMemory[12][29] ),
    .A1(net260),
    .S(net127),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(\dataMemory[12][30] ),
    .A1(net239),
    .S(net127),
    .X(_0973_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(\dataMemory[12][31] ),
    .A1(net236),
    .S(net127),
    .X(_0974_));
 sky130_fd_sc_hd__nand2_2 _3672_ (.A(_1799_),
    .B(_1810_),
    .Y(_1844_));
 sky130_fd_sc_hd__mux2_1 _3673_ (.A0(net202),
    .A1(\dataMemory[13][0] ),
    .S(net72),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _3674_ (.A0(net299),
    .A1(\dataMemory[13][1] ),
    .S(net72),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _3675_ (.A0(net258),
    .A1(\dataMemory[13][2] ),
    .S(net72),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _3676_ (.A0(net235),
    .A1(\dataMemory[13][3] ),
    .S(net72),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(net233),
    .A1(\dataMemory[13][4] ),
    .S(net72),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(net230),
    .A1(\dataMemory[13][5] ),
    .S(net72),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(net228),
    .A1(\dataMemory[13][6] ),
    .S(net72),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(net227),
    .A1(\dataMemory[13][7] ),
    .S(net73),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(net225),
    .A1(\dataMemory[13][8] ),
    .S(net72),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(net222),
    .A1(\dataMemory[13][9] ),
    .S(net72),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _3683_ (.A0(net200),
    .A1(\dataMemory[13][10] ),
    .S(net72),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _3684_ (.A0(net198),
    .A1(\dataMemory[13][11] ),
    .S(_1844_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _3685_ (.A0(net314),
    .A1(\dataMemory[13][12] ),
    .S(net72),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _3686_ (.A0(net313),
    .A1(\dataMemory[13][13] ),
    .S(net72),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _3687_ (.A0(net311),
    .A1(\dataMemory[13][14] ),
    .S(net72),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _3688_ (.A0(net309),
    .A1(\dataMemory[13][15] ),
    .S(net73),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(net307),
    .A1(\dataMemory[13][16] ),
    .S(net73),
    .X(_0991_));
 sky130_fd_sc_hd__mux2_1 _3690_ (.A0(net305),
    .A1(\dataMemory[13][17] ),
    .S(net73),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _3691_ (.A0(net302),
    .A1(\dataMemory[13][18] ),
    .S(net73),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(net300),
    .A1(\dataMemory[13][19] ),
    .S(net72),
    .X(_0994_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(net296),
    .A1(\dataMemory[13][20] ),
    .S(net72),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _3694_ (.A0(net276),
    .A1(\dataMemory[13][21] ),
    .S(net73),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _3695_ (.A0(net275),
    .A1(\dataMemory[13][22] ),
    .S(net73),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _3696_ (.A0(net22),
    .A1(\dataMemory[13][23] ),
    .S(net73),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _3697_ (.A0(net271),
    .A1(\dataMemory[13][24] ),
    .S(net73),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_1 _3698_ (.A0(net268),
    .A1(\dataMemory[13][25] ),
    .S(net73),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _3699_ (.A0(net267),
    .A1(\dataMemory[13][26] ),
    .S(net72),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _3700_ (.A0(net264),
    .A1(\dataMemory[13][27] ),
    .S(net73),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _3701_ (.A0(net262),
    .A1(\dataMemory[13][28] ),
    .S(net73),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(net261),
    .A1(\dataMemory[13][29] ),
    .S(net73),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(net239),
    .A1(\dataMemory[13][30] ),
    .S(net73),
    .X(_1005_));
 sky130_fd_sc_hd__mux2_1 _3704_ (.A0(net236),
    .A1(\dataMemory[13][31] ),
    .S(net73),
    .X(_1006_));
 sky130_fd_sc_hd__mux2_1 _3705_ (.A0(net7),
    .A1(\dataMemory[14][0] ),
    .S(net124),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(net299),
    .A1(\dataMemory[14][1] ),
    .S(net124),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _3707_ (.A0(net258),
    .A1(\dataMemory[14][2] ),
    .S(net124),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _3708_ (.A0(net235),
    .A1(\dataMemory[14][3] ),
    .S(net124),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _3709_ (.A0(net233),
    .A1(\dataMemory[14][4] ),
    .S(net124),
    .X(_1011_));
 sky130_fd_sc_hd__mux2_1 _3710_ (.A0(net230),
    .A1(\dataMemory[14][5] ),
    .S(net124),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(net228),
    .A1(\dataMemory[14][6] ),
    .S(net125),
    .X(_1013_));
 sky130_fd_sc_hd__mux2_1 _3712_ (.A0(net226),
    .A1(\dataMemory[14][7] ),
    .S(net124),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(net225),
    .A1(\dataMemory[14][8] ),
    .S(net124),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_1 _3714_ (.A0(net222),
    .A1(\dataMemory[14][9] ),
    .S(net124),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _3715_ (.A0(net200),
    .A1(\dataMemory[14][10] ),
    .S(net124),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _3716_ (.A0(net198),
    .A1(\dataMemory[14][11] ),
    .S(net125),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _3717_ (.A0(net314),
    .A1(\dataMemory[14][12] ),
    .S(net124),
    .X(_1019_));
 sky130_fd_sc_hd__mux2_1 _3718_ (.A0(net313),
    .A1(\dataMemory[14][13] ),
    .S(net124),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _3719_ (.A0(net311),
    .A1(\dataMemory[14][14] ),
    .S(net124),
    .X(_1021_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(net309),
    .A1(\dataMemory[14][15] ),
    .S(net125),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _3721_ (.A0(net307),
    .A1(\dataMemory[14][16] ),
    .S(net125),
    .X(_1023_));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(net371),
    .D(_0000_),
    .Q(\dataMemory[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(net361),
    .D(_0001_),
    .Q(\dataMemory[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(net342),
    .D(_0002_),
    .Q(\dataMemory[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(net346),
    .D(_0003_),
    .Q(\dataMemory[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(net358),
    .D(_0004_),
    .Q(\dataMemory[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(net371),
    .D(_0005_),
    .Q(\dataMemory[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(net374),
    .D(_0006_),
    .Q(\dataMemory[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(net374),
    .D(_0007_),
    .Q(\dataMemory[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(net366),
    .D(_0008_),
    .Q(\dataMemory[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(net347),
    .D(_0009_),
    .Q(\dataMemory[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(net362),
    .D(_0010_),
    .Q(\dataMemory[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(net380),
    .D(_0011_),
    .Q(\dataMemory[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(net381),
    .D(_0012_),
    .Q(\dataMemory[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(net381),
    .D(_0013_),
    .Q(\dataMemory[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(net381),
    .D(_0014_),
    .Q(\dataMemory[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(net320),
    .D(_0015_),
    .Q(\dataMemory[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(net323),
    .D(_0016_),
    .Q(\dataMemory[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(net320),
    .D(_0017_),
    .Q(\dataMemory[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(net320),
    .D(_0018_),
    .Q(\dataMemory[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(net333),
    .D(_0019_),
    .Q(\dataMemory[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(net328),
    .D(_0020_),
    .Q(\dataMemory[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(net334),
    .D(_0021_),
    .Q(\dataMemory[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(net337),
    .D(_0022_),
    .Q(\dataMemory[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(net343),
    .D(_0023_),
    .Q(\dataMemory[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(net328),
    .D(_0024_),
    .Q(\dataMemory[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(net339),
    .D(_0025_),
    .Q(\dataMemory[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(net357),
    .D(_0026_),
    .Q(\dataMemory[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(net352),
    .D(_0027_),
    .Q(\dataMemory[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(net342),
    .D(_0028_),
    .Q(\dataMemory[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(net330),
    .D(_0029_),
    .Q(\dataMemory[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(net354),
    .D(_0030_),
    .Q(\dataMemory[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(net375),
    .D(_0031_),
    .Q(\dataMemory[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(net372),
    .D(_0032_),
    .Q(\dataMemory[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(net361),
    .D(_0033_),
    .Q(\dataMemory[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(net342),
    .D(_0034_),
    .Q(\dataMemory[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(net346),
    .D(_0035_),
    .Q(\dataMemory[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(net358),
    .D(_0036_),
    .Q(\dataMemory[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(net372),
    .D(_0037_),
    .Q(\dataMemory[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(net378),
    .D(_0038_),
    .Q(\dataMemory[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(net378),
    .D(_0039_),
    .Q(\dataMemory[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(net366),
    .D(_0040_),
    .Q(\dataMemory[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(net347),
    .D(_0041_),
    .Q(\dataMemory[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(net362),
    .D(_0042_),
    .Q(\dataMemory[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(net380),
    .D(_0043_),
    .Q(\dataMemory[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(net381),
    .D(_0044_),
    .Q(\dataMemory[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(net381),
    .D(_0045_),
    .Q(\dataMemory[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(net381),
    .D(_0046_),
    .Q(\dataMemory[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(net316),
    .D(_0047_),
    .Q(\dataMemory[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(net319),
    .D(_0048_),
    .Q(\dataMemory[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(net316),
    .D(_0049_),
    .Q(\dataMemory[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3772_ (.CLK(net319),
    .D(_0050_),
    .Q(\dataMemory[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3773_ (.CLK(net334),
    .D(_0051_),
    .Q(\dataMemory[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3774_ (.CLK(net326),
    .D(_0052_),
    .Q(\dataMemory[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3775_ (.CLK(net339),
    .D(_0053_),
    .Q(\dataMemory[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3776_ (.CLK(net339),
    .D(_0054_),
    .Q(\dataMemory[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3777_ (.CLK(net328),
    .D(_0055_),
    .Q(\dataMemory[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3778_ (.CLK(net327),
    .D(_0056_),
    .Q(\dataMemory[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3779_ (.CLK(net347),
    .D(_0057_),
    .Q(\dataMemory[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3780_ (.CLK(net356),
    .D(_0058_),
    .Q(\dataMemory[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3781_ (.CLK(net355),
    .D(_0059_),
    .Q(\dataMemory[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3782_ (.CLK(net331),
    .D(_0060_),
    .Q(\dataMemory[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3783_ (.CLK(net344),
    .D(_0061_),
    .Q(\dataMemory[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3784_ (.CLK(net366),
    .D(_0062_),
    .Q(\dataMemory[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3785_ (.CLK(net356),
    .D(_0063_),
    .Q(\dataMemory[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3786_ (.CLK(net359),
    .D(_0064_),
    .Q(\dataMemory[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3787_ (.CLK(net364),
    .D(_0065_),
    .Q(\dataMemory[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3788_ (.CLK(net345),
    .D(_0066_),
    .Q(\dataMemory[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3789_ (.CLK(net349),
    .D(_0067_),
    .Q(\dataMemory[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3790_ (.CLK(net367),
    .D(_0068_),
    .Q(\dataMemory[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3791_ (.CLK(net372),
    .D(_0069_),
    .Q(\dataMemory[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3792_ (.CLK(net374),
    .D(_0070_),
    .Q(\dataMemory[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3793_ (.CLK(net381),
    .D(_0071_),
    .Q(\dataMemory[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3794_ (.CLK(net369),
    .D(_0072_),
    .Q(\dataMemory[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3795_ (.CLK(net363),
    .D(_0073_),
    .Q(\dataMemory[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3796_ (.CLK(net368),
    .D(_0074_),
    .Q(\dataMemory[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3797_ (.CLK(net383),
    .D(_0075_),
    .Q(\dataMemory[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3798_ (.CLK(net387),
    .D(_0076_),
    .Q(\dataMemory[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3799_ (.CLK(net388),
    .D(_0077_),
    .Q(\dataMemory[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3800_ (.CLK(net388),
    .D(_0078_),
    .Q(\dataMemory[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3801_ (.CLK(net316),
    .D(_0079_),
    .Q(\dataMemory[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3802_ (.CLK(net319),
    .D(_0080_),
    .Q(\dataMemory[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3803_ (.CLK(net316),
    .D(_0081_),
    .Q(\dataMemory[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3804_ (.CLK(net319),
    .D(_0082_),
    .Q(\dataMemory[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3805_ (.CLK(net335),
    .D(_0083_),
    .Q(\dataMemory[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3806_ (.CLK(net328),
    .D(_0084_),
    .Q(\dataMemory[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3807_ (.CLK(net339),
    .D(_0085_),
    .Q(\dataMemory[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3808_ (.CLK(net339),
    .D(_0086_),
    .Q(\dataMemory[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3809_ (.CLK(net326),
    .D(_0087_),
    .Q(\dataMemory[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3810_ (.CLK(net330),
    .D(_0088_),
    .Q(\dataMemory[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3811_ (.CLK(net347),
    .D(_0089_),
    .Q(\dataMemory[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3812_ (.CLK(net353),
    .D(_0090_),
    .Q(\dataMemory[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3813_ (.CLK(net352),
    .D(_0091_),
    .Q(\dataMemory[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3814_ (.CLK(net331),
    .D(_0092_),
    .Q(\dataMemory[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3815_ (.CLK(net344),
    .D(_0093_),
    .Q(\dataMemory[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3816_ (.CLK(net362),
    .D(_0094_),
    .Q(\dataMemory[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3817_ (.CLK(net356),
    .D(_0095_),
    .Q(\dataMemory[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3818_ (.CLK(net359),
    .D(_0096_),
    .Q(\dataMemory[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3819_ (.CLK(net363),
    .D(_0097_),
    .Q(\dataMemory[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3820_ (.CLK(net345),
    .D(_0098_),
    .Q(\dataMemory[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3821_ (.CLK(net348),
    .D(_0099_),
    .Q(\dataMemory[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3822_ (.CLK(net367),
    .D(_0100_),
    .Q(\dataMemory[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3823_ (.CLK(net372),
    .D(_0101_),
    .Q(\dataMemory[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3824_ (.CLK(net374),
    .D(_0102_),
    .Q(\dataMemory[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3825_ (.CLK(net381),
    .D(_0103_),
    .Q(\dataMemory[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3826_ (.CLK(net369),
    .D(_0104_),
    .Q(\dataMemory[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3827_ (.CLK(net363),
    .D(_0105_),
    .Q(\dataMemory[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3828_ (.CLK(net368),
    .D(_0106_),
    .Q(\dataMemory[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3829_ (.CLK(net383),
    .D(_0107_),
    .Q(\dataMemory[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3830_ (.CLK(net388),
    .D(_0108_),
    .Q(\dataMemory[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3831_ (.CLK(net388),
    .D(_0109_),
    .Q(\dataMemory[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3832_ (.CLK(net388),
    .D(_0110_),
    .Q(\dataMemory[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3833_ (.CLK(net316),
    .D(_0111_),
    .Q(\dataMemory[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3834_ (.CLK(net319),
    .D(_0112_),
    .Q(\dataMemory[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3835_ (.CLK(net316),
    .D(_0113_),
    .Q(\dataMemory[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3836_ (.CLK(net319),
    .D(_0114_),
    .Q(\dataMemory[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3837_ (.CLK(net335),
    .D(_0115_),
    .Q(\dataMemory[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3838_ (.CLK(net328),
    .D(_0116_),
    .Q(\dataMemory[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3839_ (.CLK(net339),
    .D(_0117_),
    .Q(\dataMemory[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3840_ (.CLK(net339),
    .D(_0118_),
    .Q(\dataMemory[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3841_ (.CLK(net328),
    .D(_0119_),
    .Q(\dataMemory[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3842_ (.CLK(net330),
    .D(_0120_),
    .Q(\dataMemory[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3843_ (.CLK(net361),
    .D(_0121_),
    .Q(\dataMemory[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3844_ (.CLK(net353),
    .D(_0122_),
    .Q(\dataMemory[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3845_ (.CLK(net353),
    .D(_0123_),
    .Q(\dataMemory[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3846_ (.CLK(net331),
    .D(_0124_),
    .Q(\dataMemory[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3847_ (.CLK(net344),
    .D(_0125_),
    .Q(\dataMemory[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3848_ (.CLK(net362),
    .D(_0126_),
    .Q(\dataMemory[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3849_ (.CLK(net356),
    .D(_0127_),
    .Q(\dataMemory[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3850_ (.CLK(net359),
    .D(_0128_),
    .Q(\dataMemory[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3851_ (.CLK(net364),
    .D(_0129_),
    .Q(\dataMemory[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3852_ (.CLK(net348),
    .D(_0130_),
    .Q(\dataMemory[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3853_ (.CLK(net349),
    .D(_0131_),
    .Q(\dataMemory[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3854_ (.CLK(net367),
    .D(_0132_),
    .Q(\dataMemory[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3855_ (.CLK(net372),
    .D(_0133_),
    .Q(\dataMemory[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3856_ (.CLK(net374),
    .D(_0134_),
    .Q(\dataMemory[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3857_ (.CLK(net381),
    .D(_0135_),
    .Q(\dataMemory[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3858_ (.CLK(net369),
    .D(_0136_),
    .Q(\dataMemory[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3859_ (.CLK(net363),
    .D(_0137_),
    .Q(\dataMemory[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3860_ (.CLK(net368),
    .D(_0138_),
    .Q(\dataMemory[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3861_ (.CLK(net383),
    .D(_0139_),
    .Q(\dataMemory[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3862_ (.CLK(net388),
    .D(_0140_),
    .Q(\dataMemory[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3863_ (.CLK(net388),
    .D(_0141_),
    .Q(\dataMemory[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3864_ (.CLK(net388),
    .D(_0142_),
    .Q(\dataMemory[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3865_ (.CLK(net321),
    .D(_0143_),
    .Q(\dataMemory[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3866_ (.CLK(net322),
    .D(_0144_),
    .Q(\dataMemory[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3867_ (.CLK(net321),
    .D(_0145_),
    .Q(\dataMemory[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3868_ (.CLK(net322),
    .D(_0146_),
    .Q(\dataMemory[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3869_ (.CLK(net334),
    .D(_0147_),
    .Q(\dataMemory[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3870_ (.CLK(net329),
    .D(_0148_),
    .Q(\dataMemory[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3871_ (.CLK(net334),
    .D(_0149_),
    .Q(\dataMemory[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3872_ (.CLK(net338),
    .D(_0150_),
    .Q(\dataMemory[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3873_ (.CLK(net335),
    .D(_0151_),
    .Q(\dataMemory[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3874_ (.CLK(net331),
    .D(_0152_),
    .Q(\dataMemory[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3875_ (.CLK(net339),
    .D(_0153_),
    .Q(\dataMemory[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3876_ (.CLK(net357),
    .D(_0154_),
    .Q(\dataMemory[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3877_ (.CLK(net352),
    .D(_0155_),
    .Q(\dataMemory[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3878_ (.CLK(net342),
    .D(_0156_),
    .Q(\dataMemory[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3879_ (.CLK(net344),
    .D(_0157_),
    .Q(\dataMemory[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3880_ (.CLK(net358),
    .D(_0158_),
    .Q(\dataMemory[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3881_ (.CLK(net376),
    .D(_0159_),
    .Q(\dataMemory[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3882_ (.CLK(net375),
    .D(_0160_),
    .Q(\dataMemory[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3883_ (.CLK(net362),
    .D(_0161_),
    .Q(\dataMemory[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3884_ (.CLK(net348),
    .D(_0162_),
    .Q(\dataMemory[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3885_ (.CLK(net349),
    .D(_0163_),
    .Q(\dataMemory[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3886_ (.CLK(net358),
    .D(_0164_),
    .Q(\dataMemory[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3887_ (.CLK(net376),
    .D(_0165_),
    .Q(\dataMemory[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3888_ (.CLK(net378),
    .D(_0166_),
    .Q(\dataMemory[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3889_ (.CLK(net378),
    .D(_0167_),
    .Q(\dataMemory[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3890_ (.CLK(net382),
    .D(_0168_),
    .Q(\dataMemory[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3891_ (.CLK(net363),
    .D(_0169_),
    .Q(\dataMemory[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3892_ (.CLK(net368),
    .D(_0170_),
    .Q(\dataMemory[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3893_ (.CLK(net381),
    .D(_0171_),
    .Q(\dataMemory[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3894_ (.CLK(net388),
    .D(_0172_),
    .Q(\dataMemory[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3895_ (.CLK(net386),
    .D(_0173_),
    .Q(\dataMemory[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3896_ (.CLK(net386),
    .D(_0174_),
    .Q(\dataMemory[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3897_ (.CLK(net316),
    .D(_0175_),
    .Q(\dataMemory[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3898_ (.CLK(net319),
    .D(_0176_),
    .Q(\dataMemory[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3899_ (.CLK(net316),
    .D(_0177_),
    .Q(\dataMemory[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3900_ (.CLK(net319),
    .D(_0178_),
    .Q(\dataMemory[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3901_ (.CLK(net334),
    .D(_0179_),
    .Q(\dataMemory[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3902_ (.CLK(net326),
    .D(_0180_),
    .Q(\dataMemory[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3903_ (.CLK(net339),
    .D(_0181_),
    .Q(\dataMemory[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3904_ (.CLK(net340),
    .D(_0182_),
    .Q(\dataMemory[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3905_ (.CLK(net326),
    .D(_0183_),
    .Q(\dataMemory[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3906_ (.CLK(net327),
    .D(_0184_),
    .Q(\dataMemory[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3907_ (.CLK(net347),
    .D(_0185_),
    .Q(\dataMemory[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3908_ (.CLK(net356),
    .D(_0186_),
    .Q(\dataMemory[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3909_ (.CLK(net354),
    .D(_0187_),
    .Q(\dataMemory[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3910_ (.CLK(net331),
    .D(_0188_),
    .Q(\dataMemory[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3911_ (.CLK(net344),
    .D(_0189_),
    .Q(\dataMemory[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3912_ (.CLK(net355),
    .D(_0190_),
    .Q(\dataMemory[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3913_ (.CLK(net356),
    .D(_0191_),
    .Q(\dataMemory[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3914_ (.CLK(net359),
    .D(_0192_),
    .Q(\dataMemory[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3915_ (.CLK(net364),
    .D(_0193_),
    .Q(\dataMemory[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3916_ (.CLK(net345),
    .D(_0194_),
    .Q(\dataMemory[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3917_ (.CLK(net348),
    .D(_0195_),
    .Q(\dataMemory[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3918_ (.CLK(net380),
    .D(_0196_),
    .Q(\dataMemory[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3919_ (.CLK(net371),
    .D(_0197_),
    .Q(\dataMemory[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3920_ (.CLK(net374),
    .D(_0198_),
    .Q(\dataMemory[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3921_ (.CLK(net374),
    .D(_0199_),
    .Q(\dataMemory[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3922_ (.CLK(net369),
    .D(_0200_),
    .Q(\dataMemory[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3923_ (.CLK(net363),
    .D(_0201_),
    .Q(\dataMemory[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3924_ (.CLK(net368),
    .D(_0202_),
    .Q(\dataMemory[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3925_ (.CLK(net382),
    .D(_0203_),
    .Q(\dataMemory[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3926_ (.CLK(net383),
    .D(_0204_),
    .Q(\dataMemory[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3927_ (.CLK(net383),
    .D(_0205_),
    .Q(\dataMemory[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3928_ (.CLK(net383),
    .D(_0206_),
    .Q(\dataMemory[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3929_ (.CLK(net316),
    .D(_0207_),
    .Q(\dataMemory[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3930_ (.CLK(net318),
    .D(_0208_),
    .Q(\dataMemory[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3931_ (.CLK(net317),
    .D(_0209_),
    .Q(\dataMemory[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3932_ (.CLK(net318),
    .D(_0210_),
    .Q(\dataMemory[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3933_ (.CLK(net333),
    .D(_0211_),
    .Q(\dataMemory[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3934_ (.CLK(net325),
    .D(_0212_),
    .Q(\dataMemory[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3935_ (.CLK(net335),
    .D(_0213_),
    .Q(\dataMemory[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3936_ (.CLK(net338),
    .D(_0214_),
    .Q(\dataMemory[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3937_ (.CLK(net325),
    .D(_0215_),
    .Q(\dataMemory[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3938_ (.CLK(net327),
    .D(_0216_),
    .Q(\dataMemory[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3939_ (.CLK(net347),
    .D(_0217_),
    .Q(\dataMemory[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3940_ (.CLK(net353),
    .D(_0218_),
    .Q(\dataMemory[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3941_ (.CLK(net354),
    .D(_0219_),
    .Q(\dataMemory[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3942_ (.CLK(net330),
    .D(_0220_),
    .Q(\dataMemory[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3943_ (.CLK(net344),
    .D(_0221_),
    .Q(\dataMemory[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3944_ (.CLK(net358),
    .D(_0222_),
    .Q(\dataMemory[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3945_ (.CLK(net356),
    .D(_0223_),
    .Q(\dataMemory[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3946_ (.CLK(net357),
    .D(_0224_),
    .Q(\dataMemory[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3947_ (.CLK(net364),
    .D(_0225_),
    .Q(\dataMemory[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3948_ (.CLK(net345),
    .D(_0226_),
    .Q(\dataMemory[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3949_ (.CLK(net348),
    .D(_0227_),
    .Q(\dataMemory[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3950_ (.CLK(net380),
    .D(_0228_),
    .Q(\dataMemory[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3951_ (.CLK(net371),
    .D(_0229_),
    .Q(\dataMemory[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3952_ (.CLK(net373),
    .D(_0230_),
    .Q(\dataMemory[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3953_ (.CLK(net373),
    .D(_0231_),
    .Q(\dataMemory[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3954_ (.CLK(net369),
    .D(_0232_),
    .Q(\dataMemory[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3955_ (.CLK(net349),
    .D(_0233_),
    .Q(\dataMemory[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3956_ (.CLK(net364),
    .D(_0234_),
    .Q(\dataMemory[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3957_ (.CLK(net382),
    .D(_0235_),
    .Q(\dataMemory[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3958_ (.CLK(net382),
    .D(_0236_),
    .Q(\dataMemory[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3959_ (.CLK(net382),
    .D(_0237_),
    .Q(\dataMemory[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3960_ (.CLK(net380),
    .D(_0238_),
    .Q(\dataMemory[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3961_ (.CLK(net316),
    .D(_0239_),
    .Q(\dataMemory[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3962_ (.CLK(net319),
    .D(_0240_),
    .Q(\dataMemory[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3963_ (.CLK(net316),
    .D(_0241_),
    .Q(\dataMemory[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3964_ (.CLK(net319),
    .D(_0242_),
    .Q(\dataMemory[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3965_ (.CLK(net333),
    .D(_0243_),
    .Q(\dataMemory[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3966_ (.CLK(net326),
    .D(_0244_),
    .Q(\dataMemory[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3967_ (.CLK(net339),
    .D(_0245_),
    .Q(\dataMemory[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3968_ (.CLK(net338),
    .D(_0246_),
    .Q(\dataMemory[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3969_ (.CLK(net326),
    .D(_0247_),
    .Q(\dataMemory[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3970_ (.CLK(net327),
    .D(_0248_),
    .Q(\dataMemory[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3971_ (.CLK(net347),
    .D(_0249_),
    .Q(\dataMemory[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3972_ (.CLK(net353),
    .D(_0250_),
    .Q(\dataMemory[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3973_ (.CLK(net354),
    .D(_0251_),
    .Q(\dataMemory[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3974_ (.CLK(net330),
    .D(_0252_),
    .Q(\dataMemory[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3975_ (.CLK(net344),
    .D(_0253_),
    .Q(\dataMemory[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3976_ (.CLK(net358),
    .D(_0254_),
    .Q(\dataMemory[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3977_ (.CLK(net356),
    .D(_0255_),
    .Q(\dataMemory[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3978_ (.CLK(net357),
    .D(_0256_),
    .Q(\dataMemory[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3979_ (.CLK(net364),
    .D(_0257_),
    .Q(\dataMemory[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3980_ (.CLK(net345),
    .D(_0258_),
    .Q(\dataMemory[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3981_ (.CLK(net348),
    .D(_0259_),
    .Q(\dataMemory[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3982_ (.CLK(net373),
    .D(_0260_),
    .Q(\dataMemory[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3983_ (.CLK(net371),
    .D(_0261_),
    .Q(\dataMemory[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3984_ (.CLK(net373),
    .D(_0262_),
    .Q(\dataMemory[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3985_ (.CLK(net373),
    .D(_0263_),
    .Q(\dataMemory[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3986_ (.CLK(net369),
    .D(_0264_),
    .Q(\dataMemory[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3987_ (.CLK(net349),
    .D(_0265_),
    .Q(\dataMemory[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3988_ (.CLK(net368),
    .D(_0266_),
    .Q(\dataMemory[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3989_ (.CLK(net382),
    .D(_0267_),
    .Q(\dataMemory[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3990_ (.CLK(net383),
    .D(_0268_),
    .Q(\dataMemory[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3991_ (.CLK(net383),
    .D(_0269_),
    .Q(\dataMemory[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3992_ (.CLK(net381),
    .D(_0270_),
    .Q(\dataMemory[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3993_ (.CLK(net317),
    .D(_0271_),
    .Q(\dataMemory[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3994_ (.CLK(net318),
    .D(_0272_),
    .Q(\dataMemory[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3995_ (.CLK(net317),
    .D(_0273_),
    .Q(\dataMemory[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3996_ (.CLK(net318),
    .D(_0274_),
    .Q(\dataMemory[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3997_ (.CLK(net333),
    .D(_0275_),
    .Q(\dataMemory[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3998_ (.CLK(net325),
    .D(_0276_),
    .Q(\dataMemory[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3999_ (.CLK(net335),
    .D(_0277_),
    .Q(\dataMemory[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4000_ (.CLK(net338),
    .D(_0278_),
    .Q(\dataMemory[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4001_ (.CLK(net325),
    .D(_0279_),
    .Q(\dataMemory[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4002_ (.CLK(net327),
    .D(_0280_),
    .Q(\dataMemory[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4003_ (.CLK(net346),
    .D(_0281_),
    .Q(\dataMemory[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4004_ (.CLK(net353),
    .D(_0282_),
    .Q(\dataMemory[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4005_ (.CLK(net354),
    .D(_0283_),
    .Q(\dataMemory[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4006_ (.CLK(net330),
    .D(_0284_),
    .Q(\dataMemory[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4007_ (.CLK(net344),
    .D(_0285_),
    .Q(\dataMemory[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4008_ (.CLK(net355),
    .D(_0286_),
    .Q(\dataMemory[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4009_ (.CLK(net356),
    .D(_0287_),
    .Q(\dataMemory[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4010_ (.CLK(net356),
    .D(_0288_),
    .Q(\dataMemory[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4011_ (.CLK(net364),
    .D(_0289_),
    .Q(\dataMemory[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4012_ (.CLK(net345),
    .D(_0290_),
    .Q(\dataMemory[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4013_ (.CLK(net348),
    .D(_0291_),
    .Q(\dataMemory[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4014_ (.CLK(net359),
    .D(_0292_),
    .Q(\dataMemory[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4015_ (.CLK(net371),
    .D(_0293_),
    .Q(\dataMemory[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4016_ (.CLK(net373),
    .D(_0294_),
    .Q(\dataMemory[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4017_ (.CLK(net373),
    .D(_0295_),
    .Q(\dataMemory[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4018_ (.CLK(net368),
    .D(_0296_),
    .Q(\dataMemory[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4019_ (.CLK(net349),
    .D(_0297_),
    .Q(\dataMemory[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4020_ (.CLK(net364),
    .D(_0298_),
    .Q(\dataMemory[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4021_ (.CLK(net382),
    .D(_0299_),
    .Q(\dataMemory[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4022_ (.CLK(net382),
    .D(_0300_),
    .Q(\dataMemory[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4023_ (.CLK(net382),
    .D(_0301_),
    .Q(\dataMemory[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4024_ (.CLK(net380),
    .D(_0302_),
    .Q(\dataMemory[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4025_ (.CLK(net316),
    .D(_0303_),
    .Q(\dataMemory[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4026_ (.CLK(net319),
    .D(_0304_),
    .Q(\dataMemory[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4027_ (.CLK(net316),
    .D(_0305_),
    .Q(\dataMemory[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4028_ (.CLK(net319),
    .D(_0306_),
    .Q(\dataMemory[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4029_ (.CLK(net336),
    .D(_0307_),
    .Q(\dataMemory[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4030_ (.CLK(net326),
    .D(_0308_),
    .Q(\dataMemory[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4031_ (.CLK(net335),
    .D(_0309_),
    .Q(\dataMemory[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4032_ (.CLK(net337),
    .D(_0310_),
    .Q(\dataMemory[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4033_ (.CLK(net326),
    .D(_0311_),
    .Q(\dataMemory[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4034_ (.CLK(net327),
    .D(_0312_),
    .Q(\dataMemory[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4035_ (.CLK(net340),
    .D(_0313_),
    .Q(\dataMemory[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4036_ (.CLK(net353),
    .D(_0314_),
    .Q(\dataMemory[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4037_ (.CLK(net354),
    .D(_0315_),
    .Q(\dataMemory[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4038_ (.CLK(net330),
    .D(_0316_),
    .Q(\dataMemory[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4039_ (.CLK(net344),
    .D(_0317_),
    .Q(\dataMemory[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4040_ (.CLK(net354),
    .D(_0318_),
    .Q(\dataMemory[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4041_ (.CLK(net357),
    .D(_0319_),
    .Q(\dataMemory[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4042_ (.CLK(net358),
    .D(_0320_),
    .Q(\dataMemory[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4043_ (.CLK(net363),
    .D(_0321_),
    .Q(\dataMemory[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4044_ (.CLK(net345),
    .D(_0322_),
    .Q(\dataMemory[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4045_ (.CLK(net348),
    .D(_0323_),
    .Q(\dataMemory[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4046_ (.CLK(net359),
    .D(_0324_),
    .Q(\dataMemory[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4047_ (.CLK(net372),
    .D(_0325_),
    .Q(\dataMemory[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4048_ (.CLK(net373),
    .D(_0326_),
    .Q(\dataMemory[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4049_ (.CLK(net374),
    .D(_0327_),
    .Q(\dataMemory[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4050_ (.CLK(net368),
    .D(_0328_),
    .Q(\dataMemory[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4051_ (.CLK(net349),
    .D(_0329_),
    .Q(\dataMemory[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4052_ (.CLK(net368),
    .D(_0330_),
    .Q(\dataMemory[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4053_ (.CLK(net382),
    .D(_0331_),
    .Q(\dataMemory[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4054_ (.CLK(net387),
    .D(_0332_),
    .Q(\dataMemory[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4055_ (.CLK(net387),
    .D(_0333_),
    .Q(\dataMemory[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4056_ (.CLK(net387),
    .D(_0334_),
    .Q(\dataMemory[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4057_ (.CLK(net317),
    .D(_0335_),
    .Q(\dataMemory[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4058_ (.CLK(net318),
    .D(_0336_),
    .Q(\dataMemory[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4059_ (.CLK(net317),
    .D(_0337_),
    .Q(\dataMemory[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4060_ (.CLK(net318),
    .D(_0338_),
    .Q(\dataMemory[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4061_ (.CLK(net322),
    .D(_0339_),
    .Q(\dataMemory[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4062_ (.CLK(net325),
    .D(_0340_),
    .Q(\dataMemory[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4063_ (.CLK(net335),
    .D(_0341_),
    .Q(\dataMemory[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4064_ (.CLK(net337),
    .D(_0342_),
    .Q(\dataMemory[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4065_ (.CLK(net325),
    .D(_0343_),
    .Q(\dataMemory[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4066_ (.CLK(net327),
    .D(_0344_),
    .Q(\dataMemory[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4067_ (.CLK(net340),
    .D(_0345_),
    .Q(\dataMemory[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4068_ (.CLK(net353),
    .D(_0346_),
    .Q(\dataMemory[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4069_ (.CLK(net340),
    .D(_0347_),
    .Q(\dataMemory[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4070_ (.CLK(net330),
    .D(_0348_),
    .Q(\dataMemory[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4071_ (.CLK(net331),
    .D(_0349_),
    .Q(\dataMemory[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4072_ (.CLK(net354),
    .D(_0350_),
    .Q(\dataMemory[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4073_ (.CLK(net356),
    .D(_0351_),
    .Q(\dataMemory[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4074_ (.CLK(net358),
    .D(_0352_),
    .Q(\dataMemory[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4075_ (.CLK(net363),
    .D(_0353_),
    .Q(\dataMemory[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4076_ (.CLK(net345),
    .D(_0354_),
    .Q(\dataMemory[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4077_ (.CLK(net348),
    .D(_0355_),
    .Q(\dataMemory[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4078_ (.CLK(net359),
    .D(_0356_),
    .Q(\dataMemory[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4079_ (.CLK(net372),
    .D(_0357_),
    .Q(\dataMemory[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4080_ (.CLK(net373),
    .D(_0358_),
    .Q(\dataMemory[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4081_ (.CLK(net374),
    .D(_0359_),
    .Q(\dataMemory[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4082_ (.CLK(net368),
    .D(_0360_),
    .Q(\dataMemory[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4083_ (.CLK(net349),
    .D(_0361_),
    .Q(\dataMemory[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4084_ (.CLK(net364),
    .D(_0362_),
    .Q(\dataMemory[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4085_ (.CLK(net382),
    .D(_0363_),
    .Q(\dataMemory[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4086_ (.CLK(net387),
    .D(_0364_),
    .Q(\dataMemory[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4087_ (.CLK(net387),
    .D(_0365_),
    .Q(\dataMemory[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4088_ (.CLK(net387),
    .D(_0366_),
    .Q(\dataMemory[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4089_ (.CLK(net316),
    .D(_0367_),
    .Q(\dataMemory[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4090_ (.CLK(net319),
    .D(_0368_),
    .Q(\dataMemory[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4091_ (.CLK(net324),
    .D(_0369_),
    .Q(\dataMemory[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4092_ (.CLK(net319),
    .D(_0370_),
    .Q(\dataMemory[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4093_ (.CLK(net333),
    .D(_0371_),
    .Q(\dataMemory[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4094_ (.CLK(net326),
    .D(_0372_),
    .Q(\dataMemory[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4095_ (.CLK(net335),
    .D(_0373_),
    .Q(\dataMemory[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4096_ (.CLK(net337),
    .D(_0374_),
    .Q(\dataMemory[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4097_ (.CLK(net326),
    .D(_0375_),
    .Q(\dataMemory[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4098_ (.CLK(net326),
    .D(_0376_),
    .Q(\dataMemory[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4099_ (.CLK(net340),
    .D(_0377_),
    .Q(\dataMemory[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4100_ (.CLK(net353),
    .D(_0378_),
    .Q(\dataMemory[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4101_ (.CLK(net354),
    .D(_0379_),
    .Q(\dataMemory[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4102_ (.CLK(net330),
    .D(_0380_),
    .Q(\dataMemory[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4103_ (.CLK(net344),
    .D(_0381_),
    .Q(\dataMemory[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4104_ (.CLK(net355),
    .D(_0382_),
    .Q(\dataMemory[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4105_ (.CLK(net356),
    .D(_0383_),
    .Q(\dataMemory[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4106_ (.CLK(net358),
    .D(_0384_),
    .Q(\dataMemory[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4107_ (.CLK(net364),
    .D(_0385_),
    .Q(\dataMemory[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4108_ (.CLK(net345),
    .D(_0386_),
    .Q(\dataMemory[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4109_ (.CLK(net348),
    .D(_0387_),
    .Q(\dataMemory[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4110_ (.CLK(net359),
    .D(_0388_),
    .Q(\dataMemory[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4111_ (.CLK(net371),
    .D(_0389_),
    .Q(\dataMemory[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4112_ (.CLK(net374),
    .D(_0390_),
    .Q(\dataMemory[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4113_ (.CLK(net374),
    .D(_0391_),
    .Q(\dataMemory[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4114_ (.CLK(net369),
    .D(_0392_),
    .Q(\dataMemory[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4115_ (.CLK(net363),
    .D(_0393_),
    .Q(\dataMemory[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4116_ (.CLK(net368),
    .D(_0394_),
    .Q(\dataMemory[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4117_ (.CLK(net382),
    .D(_0395_),
    .Q(\dataMemory[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4118_ (.CLK(net387),
    .D(_0396_),
    .Q(\dataMemory[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4119_ (.CLK(net387),
    .D(_0397_),
    .Q(\dataMemory[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4120_ (.CLK(net387),
    .D(_0398_),
    .Q(\dataMemory[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4121_ (.CLK(net317),
    .D(_0399_),
    .Q(\dataMemory[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4122_ (.CLK(net318),
    .D(_0400_),
    .Q(\dataMemory[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4123_ (.CLK(net317),
    .D(_0401_),
    .Q(\dataMemory[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4124_ (.CLK(net318),
    .D(_0402_),
    .Q(\dataMemory[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4125_ (.CLK(net321),
    .D(_0403_),
    .Q(\dataMemory[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4126_ (.CLK(net325),
    .D(_0404_),
    .Q(\dataMemory[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4127_ (.CLK(net336),
    .D(_0405_),
    .Q(\dataMemory[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4128_ (.CLK(net337),
    .D(_0406_),
    .Q(\dataMemory[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4129_ (.CLK(net325),
    .D(_0407_),
    .Q(\dataMemory[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4130_ (.CLK(net327),
    .D(_0408_),
    .Q(\dataMemory[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4131_ (.CLK(net339),
    .D(_0409_),
    .Q(\dataMemory[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4132_ (.CLK(net353),
    .D(_0410_),
    .Q(\dataMemory[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4133_ (.CLK(net340),
    .D(_0411_),
    .Q(\dataMemory[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4134_ (.CLK(net330),
    .D(_0412_),
    .Q(\dataMemory[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4135_ (.CLK(net331),
    .D(_0413_),
    .Q(\dataMemory[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4136_ (.CLK(net354),
    .D(_0414_),
    .Q(\dataMemory[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4137_ (.CLK(net356),
    .D(_0415_),
    .Q(\dataMemory[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4138_ (.CLK(net358),
    .D(_0416_),
    .Q(\dataMemory[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4139_ (.CLK(net363),
    .D(_0417_),
    .Q(\dataMemory[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4140_ (.CLK(net345),
    .D(_0418_),
    .Q(\dataMemory[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4141_ (.CLK(net348),
    .D(_0419_),
    .Q(\dataMemory[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4142_ (.CLK(net358),
    .D(_0420_),
    .Q(\dataMemory[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4143_ (.CLK(net372),
    .D(_0421_),
    .Q(\dataMemory[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4144_ (.CLK(net373),
    .D(_0422_),
    .Q(\dataMemory[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4145_ (.CLK(net374),
    .D(_0423_),
    .Q(\dataMemory[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4146_ (.CLK(net368),
    .D(_0424_),
    .Q(\dataMemory[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4147_ (.CLK(net349),
    .D(_0425_),
    .Q(\dataMemory[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4148_ (.CLK(net364),
    .D(_0426_),
    .Q(\dataMemory[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4149_ (.CLK(net382),
    .D(_0427_),
    .Q(\dataMemory[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4150_ (.CLK(net387),
    .D(_0428_),
    .Q(\dataMemory[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4151_ (.CLK(net387),
    .D(_0429_),
    .Q(\dataMemory[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4152_ (.CLK(net387),
    .D(_0430_),
    .Q(\dataMemory[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4153_ (.CLK(net317),
    .D(_0431_),
    .Q(\dataMemory[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4154_ (.CLK(net318),
    .D(_0432_),
    .Q(\dataMemory[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4155_ (.CLK(net317),
    .D(_0433_),
    .Q(\dataMemory[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4156_ (.CLK(net318),
    .D(_0434_),
    .Q(\dataMemory[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4157_ (.CLK(net336),
    .D(_0435_),
    .Q(\dataMemory[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4158_ (.CLK(net325),
    .D(_0436_),
    .Q(\dataMemory[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4159_ (.CLK(net335),
    .D(_0437_),
    .Q(\dataMemory[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4160_ (.CLK(net337),
    .D(_0438_),
    .Q(\dataMemory[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4161_ (.CLK(net325),
    .D(_0439_),
    .Q(\dataMemory[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4162_ (.CLK(net327),
    .D(_0440_),
    .Q(\dataMemory[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4163_ (.CLK(net346),
    .D(_0441_),
    .Q(\dataMemory[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4164_ (.CLK(net356),
    .D(_0442_),
    .Q(\dataMemory[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4165_ (.CLK(net352),
    .D(_0443_),
    .Q(\dataMemory[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4166_ (.CLK(net330),
    .D(_0444_),
    .Q(\dataMemory[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4167_ (.CLK(net344),
    .D(_0445_),
    .Q(\dataMemory[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4168_ (.CLK(net361),
    .D(_0446_),
    .Q(\dataMemory[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4169_ (.CLK(net356),
    .D(_0447_),
    .Q(\dataMemory[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4170_ (.CLK(net357),
    .D(_0448_),
    .Q(\dataMemory[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4171_ (.CLK(net364),
    .D(_0449_),
    .Q(\dataMemory[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4172_ (.CLK(net345),
    .D(_0450_),
    .Q(\dataMemory[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4173_ (.CLK(net348),
    .D(_0451_),
    .Q(\dataMemory[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4174_ (.CLK(net366),
    .D(_0452_),
    .Q(\dataMemory[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4175_ (.CLK(net371),
    .D(_0453_),
    .Q(\dataMemory[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4176_ (.CLK(net373),
    .D(_0454_),
    .Q(\dataMemory[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4177_ (.CLK(net381),
    .D(_0455_),
    .Q(\dataMemory[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4178_ (.CLK(net369),
    .D(_0456_),
    .Q(\dataMemory[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4179_ (.CLK(net363),
    .D(_0457_),
    .Q(\dataMemory[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4180_ (.CLK(net368),
    .D(_0458_),
    .Q(\dataMemory[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4181_ (.CLK(net382),
    .D(_0459_),
    .Q(\dataMemory[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4182_ (.CLK(net387),
    .D(_0460_),
    .Q(\dataMemory[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4183_ (.CLK(net387),
    .D(_0461_),
    .Q(\dataMemory[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4184_ (.CLK(net383),
    .D(_0462_),
    .Q(\dataMemory[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4185_ (.CLK(net321),
    .D(_0463_),
    .Q(\dataMemory[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4186_ (.CLK(net322),
    .D(_0464_),
    .Q(\dataMemory[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4187_ (.CLK(net321),
    .D(_0465_),
    .Q(\dataMemory[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4188_ (.CLK(net322),
    .D(_0466_),
    .Q(\dataMemory[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4189_ (.CLK(net334),
    .D(_0467_),
    .Q(\dataMemory[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4190_ (.CLK(net329),
    .D(_0468_),
    .Q(\dataMemory[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4191_ (.CLK(net337),
    .D(_0469_),
    .Q(\dataMemory[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4192_ (.CLK(net338),
    .D(_0470_),
    .Q(\dataMemory[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4193_ (.CLK(net335),
    .D(_0471_),
    .Q(\dataMemory[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4194_ (.CLK(net331),
    .D(_0472_),
    .Q(\dataMemory[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4195_ (.CLK(net354),
    .D(_0473_),
    .Q(\dataMemory[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4196_ (.CLK(net357),
    .D(_0474_),
    .Q(\dataMemory[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4197_ (.CLK(net352),
    .D(_0475_),
    .Q(\dataMemory[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4198_ (.CLK(net342),
    .D(_0476_),
    .Q(\dataMemory[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4199_ (.CLK(net344),
    .D(_0477_),
    .Q(\dataMemory[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4200_ (.CLK(net358),
    .D(_0478_),
    .Q(\dataMemory[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4201_ (.CLK(net376),
    .D(_0479_),
    .Q(\dataMemory[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4202_ (.CLK(net375),
    .D(_0480_),
    .Q(\dataMemory[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4203_ (.CLK(net362),
    .D(_0481_),
    .Q(\dataMemory[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4204_ (.CLK(net348),
    .D(_0482_),
    .Q(\dataMemory[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4205_ (.CLK(net349),
    .D(_0483_),
    .Q(\dataMemory[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4206_ (.CLK(net359),
    .D(_0484_),
    .Q(\dataMemory[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4207_ (.CLK(net376),
    .D(_0485_),
    .Q(\dataMemory[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4208_ (.CLK(net379),
    .D(_0486_),
    .Q(\dataMemory[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4209_ (.CLK(net379),
    .D(_0487_),
    .Q(\dataMemory[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4210_ (.CLK(net382),
    .D(_0488_),
    .Q(\dataMemory[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4211_ (.CLK(net363),
    .D(_0489_),
    .Q(\dataMemory[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4212_ (.CLK(net368),
    .D(_0490_),
    .Q(\dataMemory[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4213_ (.CLK(net381),
    .D(_0491_),
    .Q(\dataMemory[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4214_ (.CLK(net388),
    .D(_0492_),
    .Q(\dataMemory[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4215_ (.CLK(net386),
    .D(_0493_),
    .Q(\dataMemory[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4216_ (.CLK(net386),
    .D(_0494_),
    .Q(\dataMemory[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4217_ (.CLK(net317),
    .D(_0495_),
    .Q(\dataMemory[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4218_ (.CLK(net318),
    .D(_0496_),
    .Q(\dataMemory[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4219_ (.CLK(net317),
    .D(_0497_),
    .Q(\dataMemory[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4220_ (.CLK(net318),
    .D(_0498_),
    .Q(\dataMemory[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4221_ (.CLK(net336),
    .D(_0499_),
    .Q(\dataMemory[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4222_ (.CLK(net325),
    .D(_0500_),
    .Q(\dataMemory[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4223_ (.CLK(net335),
    .D(_0501_),
    .Q(\dataMemory[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4224_ (.CLK(net338),
    .D(_0502_),
    .Q(\dataMemory[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4225_ (.CLK(net325),
    .D(_0503_),
    .Q(\dataMemory[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4226_ (.CLK(net327),
    .D(_0504_),
    .Q(\dataMemory[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4227_ (.CLK(net346),
    .D(_0505_),
    .Q(\dataMemory[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4228_ (.CLK(net353),
    .D(_0506_),
    .Q(\dataMemory[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4229_ (.CLK(net338),
    .D(_0507_),
    .Q(\dataMemory[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4230_ (.CLK(net330),
    .D(_0508_),
    .Q(\dataMemory[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4231_ (.CLK(net331),
    .D(_0509_),
    .Q(\dataMemory[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4232_ (.CLK(net361),
    .D(_0510_),
    .Q(\dataMemory[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4233_ (.CLK(net357),
    .D(_0511_),
    .Q(\dataMemory[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4234_ (.CLK(net358),
    .D(_0512_),
    .Q(\dataMemory[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4235_ (.CLK(net363),
    .D(_0513_),
    .Q(\dataMemory[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4236_ (.CLK(net344),
    .D(_0514_),
    .Q(\dataMemory[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4237_ (.CLK(net349),
    .D(_0515_),
    .Q(\dataMemory[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4238_ (.CLK(net366),
    .D(_0516_),
    .Q(\dataMemory[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4239_ (.CLK(net357),
    .D(_0517_),
    .Q(\dataMemory[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4240_ (.CLK(net373),
    .D(_0518_),
    .Q(\dataMemory[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4241_ (.CLK(net380),
    .D(_0519_),
    .Q(\dataMemory[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4242_ (.CLK(net369),
    .D(_0520_),
    .Q(\dataMemory[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4243_ (.CLK(net349),
    .D(_0521_),
    .Q(\dataMemory[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4244_ (.CLK(net364),
    .D(_0522_),
    .Q(\dataMemory[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4245_ (.CLK(net382),
    .D(_0523_),
    .Q(\dataMemory[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4246_ (.CLK(net383),
    .D(_0524_),
    .Q(\dataMemory[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4247_ (.CLK(net383),
    .D(_0525_),
    .Q(\dataMemory[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4248_ (.CLK(net383),
    .D(_0526_),
    .Q(\dataMemory[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4249_ (.CLK(net320),
    .D(_0527_),
    .Q(\dataMemory[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4250_ (.CLK(net323),
    .D(_0528_),
    .Q(\dataMemory[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4251_ (.CLK(net320),
    .D(_0529_),
    .Q(\dataMemory[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4252_ (.CLK(net323),
    .D(_0530_),
    .Q(\dataMemory[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4253_ (.CLK(net333),
    .D(_0531_),
    .Q(\dataMemory[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4254_ (.CLK(net328),
    .D(_0532_),
    .Q(\dataMemory[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4255_ (.CLK(net334),
    .D(_0533_),
    .Q(\dataMemory[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4256_ (.CLK(net337),
    .D(_0534_),
    .Q(\dataMemory[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4257_ (.CLK(net336),
    .D(_0535_),
    .Q(\dataMemory[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4258_ (.CLK(net328),
    .D(_0536_),
    .Q(\dataMemory[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4259_ (.CLK(net340),
    .D(_0537_),
    .Q(\dataMemory[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4260_ (.CLK(net357),
    .D(_0538_),
    .Q(\dataMemory[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4261_ (.CLK(net352),
    .D(_0539_),
    .Q(\dataMemory[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4262_ (.CLK(net343),
    .D(_0540_),
    .Q(\dataMemory[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4263_ (.CLK(net329),
    .D(_0541_),
    .Q(\dataMemory[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4264_ (.CLK(net355),
    .D(_0542_),
    .Q(\dataMemory[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4265_ (.CLK(net375),
    .D(_0543_),
    .Q(\dataMemory[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4266_ (.CLK(net372),
    .D(_0544_),
    .Q(\dataMemory[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4267_ (.CLK(net361),
    .D(_0545_),
    .Q(\dataMemory[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4268_ (.CLK(net342),
    .D(_0546_),
    .Q(\dataMemory[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4269_ (.CLK(net346),
    .D(_0547_),
    .Q(\dataMemory[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4270_ (.CLK(net359),
    .D(_0548_),
    .Q(\dataMemory[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4271_ (.CLK(net375),
    .D(_0549_),
    .Q(\dataMemory[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4272_ (.CLK(net378),
    .D(_0550_),
    .Q(\dataMemory[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4273_ (.CLK(net378),
    .D(_0551_),
    .Q(\dataMemory[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4274_ (.CLK(net367),
    .D(_0552_),
    .Q(\dataMemory[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4275_ (.CLK(net347),
    .D(_0553_),
    .Q(\dataMemory[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4276_ (.CLK(net362),
    .D(_0554_),
    .Q(\dataMemory[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4277_ (.CLK(net380),
    .D(_0555_),
    .Q(\dataMemory[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4278_ (.CLK(net385),
    .D(_0556_),
    .Q(\dataMemory[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4279_ (.CLK(net385),
    .D(_0557_),
    .Q(\dataMemory[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4280_ (.CLK(net385),
    .D(_0558_),
    .Q(\dataMemory[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4281_ (.CLK(net333),
    .D(_0559_),
    .Q(\dataMemory[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4282_ (.CLK(net322),
    .D(_0560_),
    .Q(\dataMemory[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4283_ (.CLK(net321),
    .D(_0561_),
    .Q(\dataMemory[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4284_ (.CLK(net322),
    .D(_0562_),
    .Q(\dataMemory[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4285_ (.CLK(net333),
    .D(_0563_),
    .Q(\dataMemory[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4286_ (.CLK(net329),
    .D(_0564_),
    .Q(\dataMemory[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4287_ (.CLK(net337),
    .D(_0565_),
    .Q(\dataMemory[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4288_ (.CLK(net338),
    .D(_0566_),
    .Q(\dataMemory[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4289_ (.CLK(net336),
    .D(_0567_),
    .Q(\dataMemory[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4290_ (.CLK(net329),
    .D(_0568_),
    .Q(\dataMemory[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4291_ (.CLK(net354),
    .D(_0569_),
    .Q(\dataMemory[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4292_ (.CLK(net371),
    .D(_0570_),
    .Q(\dataMemory[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4293_ (.CLK(net352),
    .D(_0571_),
    .Q(\dataMemory[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4294_ (.CLK(net342),
    .D(_0572_),
    .Q(\dataMemory[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4295_ (.CLK(net343),
    .D(_0573_),
    .Q(\dataMemory[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4296_ (.CLK(net355),
    .D(_0574_),
    .Q(\dataMemory[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4297_ (.CLK(net376),
    .D(_0575_),
    .Q(\dataMemory[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4298_ (.CLK(net376),
    .D(_0576_),
    .Q(\dataMemory[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4299_ (.CLK(net362),
    .D(_0577_),
    .Q(\dataMemory[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4300_ (.CLK(net342),
    .D(_0578_),
    .Q(\dataMemory[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4301_ (.CLK(net347),
    .D(_0579_),
    .Q(\dataMemory[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4302_ (.CLK(net359),
    .D(_0580_),
    .Q(\dataMemory[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4303_ (.CLK(net376),
    .D(_0581_),
    .Q(\dataMemory[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4304_ (.CLK(net379),
    .D(_0582_),
    .Q(\dataMemory[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4305_ (.CLK(net379),
    .D(_0583_),
    .Q(\dataMemory[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4306_ (.CLK(net367),
    .D(_0584_),
    .Q(\dataMemory[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4307_ (.CLK(net361),
    .D(_0585_),
    .Q(\dataMemory[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4308_ (.CLK(net366),
    .D(_0586_),
    .Q(\dataMemory[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4309_ (.CLK(net380),
    .D(_0587_),
    .Q(\dataMemory[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4310_ (.CLK(net386),
    .D(_0588_),
    .Q(\dataMemory[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4311_ (.CLK(net386),
    .D(_0589_),
    .Q(\dataMemory[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4312_ (.CLK(net386),
    .D(_0590_),
    .Q(\dataMemory[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4313_ (.CLK(net333),
    .D(_0591_),
    .Q(\dataMemory[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4314_ (.CLK(net323),
    .D(_0592_),
    .Q(\dataMemory[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4315_ (.CLK(net321),
    .D(_0593_),
    .Q(\dataMemory[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4316_ (.CLK(net322),
    .D(_0594_),
    .Q(\dataMemory[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4317_ (.CLK(net334),
    .D(_0595_),
    .Q(\dataMemory[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4318_ (.CLK(net329),
    .D(_0596_),
    .Q(\dataMemory[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4319_ (.CLK(net337),
    .D(_0597_),
    .Q(\dataMemory[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4320_ (.CLK(net338),
    .D(_0598_),
    .Q(\dataMemory[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4321_ (.CLK(net336),
    .D(_0599_),
    .Q(\dataMemory[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4322_ (.CLK(net329),
    .D(_0600_),
    .Q(\dataMemory[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4323_ (.CLK(net340),
    .D(_0601_),
    .Q(\dataMemory[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4324_ (.CLK(net371),
    .D(_0602_),
    .Q(\dataMemory[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4325_ (.CLK(net352),
    .D(_0603_),
    .Q(\dataMemory[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4326_ (.CLK(net342),
    .D(_0604_),
    .Q(\dataMemory[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4327_ (.CLK(net343),
    .D(_0605_),
    .Q(\dataMemory[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4328_ (.CLK(net355),
    .D(_0606_),
    .Q(\dataMemory[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4329_ (.CLK(net376),
    .D(_0607_),
    .Q(\dataMemory[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4330_ (.CLK(net376),
    .D(_0608_),
    .Q(\dataMemory[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4331_ (.CLK(net362),
    .D(_0609_),
    .Q(\dataMemory[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4332_ (.CLK(net346),
    .D(_0610_),
    .Q(\dataMemory[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4333_ (.CLK(net347),
    .D(_0611_),
    .Q(\dataMemory[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4334_ (.CLK(net359),
    .D(_0612_),
    .Q(\dataMemory[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4335_ (.CLK(net376),
    .D(_0613_),
    .Q(\dataMemory[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4336_ (.CLK(net379),
    .D(_0614_),
    .Q(\dataMemory[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4337_ (.CLK(net379),
    .D(_0615_),
    .Q(\dataMemory[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4338_ (.CLK(net367),
    .D(_0616_),
    .Q(\dataMemory[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4339_ (.CLK(net361),
    .D(_0617_),
    .Q(\dataMemory[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4340_ (.CLK(net366),
    .D(_0618_),
    .Q(\dataMemory[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4341_ (.CLK(net380),
    .D(_0619_),
    .Q(\dataMemory[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4342_ (.CLK(net386),
    .D(_0620_),
    .Q(\dataMemory[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4343_ (.CLK(net386),
    .D(_0621_),
    .Q(\dataMemory[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4344_ (.CLK(net385),
    .D(_0622_),
    .Q(\dataMemory[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4345_ (.CLK(net321),
    .D(_0623_),
    .Q(\dataMemory[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4346_ (.CLK(net322),
    .D(_0624_),
    .Q(\dataMemory[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4347_ (.CLK(net321),
    .D(_0625_),
    .Q(\dataMemory[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4348_ (.CLK(net322),
    .D(_0626_),
    .Q(\dataMemory[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4349_ (.CLK(net334),
    .D(_0627_),
    .Q(\dataMemory[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4350_ (.CLK(net322),
    .D(_0628_),
    .Q(\dataMemory[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4351_ (.CLK(net341),
    .D(_0629_),
    .Q(\dataMemory[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4352_ (.CLK(net338),
    .D(_0630_),
    .Q(\dataMemory[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4353_ (.CLK(net335),
    .D(_0631_),
    .Q(\dataMemory[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4354_ (.CLK(net331),
    .D(_0632_),
    .Q(\dataMemory[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4355_ (.CLK(net340),
    .D(_0633_),
    .Q(\dataMemory[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4356_ (.CLK(net357),
    .D(_0634_),
    .Q(\dataMemory[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4357_ (.CLK(net352),
    .D(_0635_),
    .Q(\dataMemory[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4358_ (.CLK(net343),
    .D(_0636_),
    .Q(\dataMemory[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4359_ (.CLK(net344),
    .D(_0637_),
    .Q(\dataMemory[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4360_ (.CLK(net355),
    .D(_0638_),
    .Q(\dataMemory[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4361_ (.CLK(net376),
    .D(_0639_),
    .Q(\dataMemory[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4362_ (.CLK(net375),
    .D(_0640_),
    .Q(\dataMemory[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4363_ (.CLK(net361),
    .D(_0641_),
    .Q(\dataMemory[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4364_ (.CLK(net345),
    .D(_0642_),
    .Q(\dataMemory[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4365_ (.CLK(net348),
    .D(_0643_),
    .Q(\dataMemory[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4366_ (.CLK(net359),
    .D(_0644_),
    .Q(\dataMemory[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4367_ (.CLK(net377),
    .D(_0645_),
    .Q(\dataMemory[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4368_ (.CLK(net379),
    .D(_0646_),
    .Q(\dataMemory[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4369_ (.CLK(net379),
    .D(_0647_),
    .Q(\dataMemory[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4370_ (.CLK(net369),
    .D(_0648_),
    .Q(\dataMemory[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4371_ (.CLK(net363),
    .D(_0649_),
    .Q(\dataMemory[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4372_ (.CLK(net368),
    .D(_0650_),
    .Q(\dataMemory[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4373_ (.CLK(net381),
    .D(_0651_),
    .Q(\dataMemory[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4374_ (.CLK(net388),
    .D(_0652_),
    .Q(\dataMemory[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4375_ (.CLK(net386),
    .D(_0653_),
    .Q(\dataMemory[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4376_ (.CLK(net386),
    .D(_0654_),
    .Q(\dataMemory[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4377_ (.CLK(net317),
    .D(_0655_),
    .Q(\dataMemory[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4378_ (.CLK(net318),
    .D(_0656_),
    .Q(\dataMemory[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4379_ (.CLK(net317),
    .D(_0657_),
    .Q(\dataMemory[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4380_ (.CLK(net318),
    .D(_0658_),
    .Q(\dataMemory[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4381_ (.CLK(net336),
    .D(_0659_),
    .Q(\dataMemory[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4382_ (.CLK(net325),
    .D(_0660_),
    .Q(\dataMemory[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4383_ (.CLK(net335),
    .D(_0661_),
    .Q(\dataMemory[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4384_ (.CLK(net338),
    .D(_0662_),
    .Q(\dataMemory[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4385_ (.CLK(net325),
    .D(_0663_),
    .Q(\dataMemory[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4386_ (.CLK(net327),
    .D(_0664_),
    .Q(\dataMemory[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4387_ (.CLK(net346),
    .D(_0665_),
    .Q(\dataMemory[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4388_ (.CLK(net353),
    .D(_0666_),
    .Q(\dataMemory[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4389_ (.CLK(net352),
    .D(_0667_),
    .Q(\dataMemory[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4390_ (.CLK(net330),
    .D(_0668_),
    .Q(\dataMemory[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4391_ (.CLK(net331),
    .D(_0669_),
    .Q(\dataMemory[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4392_ (.CLK(net361),
    .D(_0670_),
    .Q(\dataMemory[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4393_ (.CLK(net357),
    .D(_0671_),
    .Q(\dataMemory[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4394_ (.CLK(net358),
    .D(_0672_),
    .Q(\dataMemory[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4395_ (.CLK(net364),
    .D(_0673_),
    .Q(\dataMemory[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4396_ (.CLK(net345),
    .D(_0674_),
    .Q(\dataMemory[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4397_ (.CLK(net349),
    .D(_0675_),
    .Q(\dataMemory[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4398_ (.CLK(net366),
    .D(_0676_),
    .Q(\dataMemory[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4399_ (.CLK(net371),
    .D(_0677_),
    .Q(\dataMemory[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4400_ (.CLK(net373),
    .D(_0678_),
    .Q(\dataMemory[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4401_ (.CLK(net380),
    .D(_0679_),
    .Q(\dataMemory[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4402_ (.CLK(net369),
    .D(_0680_),
    .Q(\dataMemory[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4403_ (.CLK(net349),
    .D(_0681_),
    .Q(\dataMemory[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4404_ (.CLK(net364),
    .D(_0682_),
    .Q(\dataMemory[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4405_ (.CLK(net384),
    .D(_0683_),
    .Q(\dataMemory[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(net383),
    .D(_0684_),
    .Q(\dataMemory[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4407_ (.CLK(net383),
    .D(_0685_),
    .Q(\dataMemory[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4408_ (.CLK(net383),
    .D(_0686_),
    .Q(\dataMemory[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4409_ (.CLK(net316),
    .D(_0687_),
    .Q(\dataMemory[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4410_ (.CLK(net319),
    .D(_0688_),
    .Q(\dataMemory[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(net324),
    .D(_0689_),
    .Q(\dataMemory[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(net319),
    .D(_0690_),
    .Q(\dataMemory[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(net335),
    .D(_0691_),
    .Q(\dataMemory[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(net326),
    .D(_0692_),
    .Q(\dataMemory[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(net335),
    .D(_0693_),
    .Q(\dataMemory[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(net339),
    .D(_0694_),
    .Q(\dataMemory[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(net326),
    .D(_0695_),
    .Q(\dataMemory[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(net330),
    .D(_0696_),
    .Q(\dataMemory[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(net347),
    .D(_0697_),
    .Q(\dataMemory[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(net353),
    .D(_0698_),
    .Q(\dataMemory[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(net352),
    .D(_0699_),
    .Q(\dataMemory[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(net330),
    .D(_0700_),
    .Q(\dataMemory[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(net351),
    .D(_0701_),
    .Q(\dataMemory[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(net362),
    .D(_0702_),
    .Q(\dataMemory[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(net356),
    .D(_0703_),
    .Q(\dataMemory[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(net357),
    .D(_0704_),
    .Q(\dataMemory[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(net363),
    .D(_0705_),
    .Q(\dataMemory[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(net345),
    .D(_0706_),
    .Q(\dataMemory[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(net350),
    .D(_0707_),
    .Q(\dataMemory[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(net367),
    .D(_0708_),
    .Q(\dataMemory[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(net372),
    .D(_0709_),
    .Q(\dataMemory[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(net374),
    .D(_0710_),
    .Q(\dataMemory[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(net374),
    .D(_0711_),
    .Q(\dataMemory[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(net369),
    .D(_0712_),
    .Q(\dataMemory[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(net365),
    .D(_0713_),
    .Q(\dataMemory[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(net369),
    .D(_0714_),
    .Q(\dataMemory[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4437_ (.CLK(net384),
    .D(_0715_),
    .Q(\dataMemory[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(net388),
    .D(_0716_),
    .Q(\dataMemory[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(net388),
    .D(_0717_),
    .Q(\dataMemory[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4440_ (.CLK(net388),
    .D(_0718_),
    .Q(\dataMemory[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(net333),
    .D(_0719_),
    .Q(\dataMemory[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4442_ (.CLK(net322),
    .D(_0720_),
    .Q(\dataMemory[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(net321),
    .D(_0721_),
    .Q(\dataMemory[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(net322),
    .D(_0722_),
    .Q(\dataMemory[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(net333),
    .D(_0723_),
    .Q(\dataMemory[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(net329),
    .D(_0724_),
    .Q(\dataMemory[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(net337),
    .D(_0725_),
    .Q(\dataMemory[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(net338),
    .D(_0726_),
    .Q(\dataMemory[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(net336),
    .D(_0727_),
    .Q(\dataMemory[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(net329),
    .D(_0728_),
    .Q(\dataMemory[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(net354),
    .D(_0729_),
    .Q(\dataMemory[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(net371),
    .D(_0730_),
    .Q(\dataMemory[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(net370),
    .D(_0731_),
    .Q(\dataMemory[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(net342),
    .D(_0732_),
    .Q(\dataMemory[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(net343),
    .D(_0733_),
    .Q(\dataMemory[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(net355),
    .D(_0734_),
    .Q(\dataMemory[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(net376),
    .D(_0735_),
    .Q(\dataMemory[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(net376),
    .D(_0736_),
    .Q(\dataMemory[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(net362),
    .D(_0737_),
    .Q(\dataMemory[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(net346),
    .D(_0738_),
    .Q(\dataMemory[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(net347),
    .D(_0739_),
    .Q(\dataMemory[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(net373),
    .D(_0740_),
    .Q(\dataMemory[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(net377),
    .D(_0741_),
    .Q(\dataMemory[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(net379),
    .D(_0742_),
    .Q(\dataMemory[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(net379),
    .D(_0743_),
    .Q(\dataMemory[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(net367),
    .D(_0744_),
    .Q(\dataMemory[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(net361),
    .D(_0745_),
    .Q(\dataMemory[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(net366),
    .D(_0746_),
    .Q(\dataMemory[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(net380),
    .D(_0747_),
    .Q(\dataMemory[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(net386),
    .D(_0748_),
    .Q(\dataMemory[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(net386),
    .D(_0749_),
    .Q(\dataMemory[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(net386),
    .D(_0750_),
    .Q(\dataMemory[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(net317),
    .D(_0751_),
    .Q(\dataMemory[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(net318),
    .D(_0752_),
    .Q(\dataMemory[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(net317),
    .D(_0753_),
    .Q(\dataMemory[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(net318),
    .D(_0754_),
    .Q(\dataMemory[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(net336),
    .D(_0755_),
    .Q(\dataMemory[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(net325),
    .D(_0756_),
    .Q(\dataMemory[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(net335),
    .D(_0757_),
    .Q(\dataMemory[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(net339),
    .D(_0758_),
    .Q(\dataMemory[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(net325),
    .D(_0759_),
    .Q(\dataMemory[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(net327),
    .D(_0760_),
    .Q(\dataMemory[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(net346),
    .D(_0761_),
    .Q(\dataMemory[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4484_ (.CLK(net370),
    .D(_0762_),
    .Q(\dataMemory[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4485_ (.CLK(net353),
    .D(_0763_),
    .Q(\dataMemory[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(net330),
    .D(_0764_),
    .Q(\dataMemory[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(net331),
    .D(_0765_),
    .Q(\dataMemory[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(net361),
    .D(_0766_),
    .Q(\dataMemory[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(net357),
    .D(_0767_),
    .Q(\dataMemory[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(net358),
    .D(_0768_),
    .Q(\dataMemory[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(net365),
    .D(_0769_),
    .Q(\dataMemory[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(net351),
    .D(_0770_),
    .Q(\dataMemory[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(net349),
    .D(_0771_),
    .Q(\dataMemory[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(net366),
    .D(_0772_),
    .Q(\dataMemory[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(net371),
    .D(_0773_),
    .Q(\dataMemory[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(net373),
    .D(_0774_),
    .Q(\dataMemory[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(net380),
    .D(_0775_),
    .Q(\dataMemory[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(net369),
    .D(_0776_),
    .Q(\dataMemory[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(net365),
    .D(_0777_),
    .Q(\dataMemory[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(net369),
    .D(_0778_),
    .Q(\dataMemory[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(net384),
    .D(_0779_),
    .Q(\dataMemory[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(net387),
    .D(_0780_),
    .Q(\dataMemory[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(net384),
    .D(_0781_),
    .Q(\dataMemory[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(net383),
    .D(_0782_),
    .Q(\dataMemory[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(net321),
    .D(_0783_),
    .Q(\dataMemory[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(net322),
    .D(_0784_),
    .Q(\dataMemory[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(net321),
    .D(_0785_),
    .Q(\dataMemory[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(net322),
    .D(_0786_),
    .Q(\dataMemory[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(net333),
    .D(_0787_),
    .Q(\dataMemory[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(net329),
    .D(_0788_),
    .Q(\dataMemory[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(net334),
    .D(_0789_),
    .Q(\dataMemory[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(net338),
    .D(_0790_),
    .Q(\dataMemory[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(net336),
    .D(_0791_),
    .Q(\dataMemory[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(net329),
    .D(_0792_),
    .Q(\dataMemory[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(net354),
    .D(_0793_),
    .Q(\dataMemory[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(net371),
    .D(_0794_),
    .Q(\dataMemory[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(net370),
    .D(_0795_),
    .Q(\dataMemory[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(net342),
    .D(_0796_),
    .Q(\dataMemory[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(net343),
    .D(_0797_),
    .Q(\dataMemory[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(net355),
    .D(_0798_),
    .Q(\dataMemory[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(net376),
    .D(_0799_),
    .Q(\dataMemory[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(net375),
    .D(_0800_),
    .Q(\dataMemory[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(net362),
    .D(_0801_),
    .Q(\dataMemory[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(net342),
    .D(_0802_),
    .Q(\dataMemory[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(net347),
    .D(_0803_),
    .Q(\dataMemory[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(net373),
    .D(_0804_),
    .Q(\dataMemory[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(net377),
    .D(_0805_),
    .Q(\dataMemory[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(net379),
    .D(_0806_),
    .Q(\dataMemory[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(net379),
    .D(_0807_),
    .Q(\dataMemory[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(net367),
    .D(_0808_),
    .Q(\dataMemory[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(net347),
    .D(_0809_),
    .Q(\dataMemory[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(net366),
    .D(_0810_),
    .Q(\dataMemory[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(net380),
    .D(_0811_),
    .Q(\dataMemory[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(net386),
    .D(_0812_),
    .Q(\dataMemory[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(net385),
    .D(_0813_),
    .Q(\dataMemory[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(net386),
    .D(_0814_),
    .Q(\dataMemory[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(net320),
    .D(_0815_),
    .Q(\dataMemory[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(net323),
    .D(_0816_),
    .Q(\dataMemory[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(net320),
    .D(_0817_),
    .Q(\dataMemory[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(net323),
    .D(_0818_),
    .Q(\dataMemory[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(net333),
    .D(_0819_),
    .Q(\dataMemory[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(net328),
    .D(_0820_),
    .Q(\dataMemory[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(net334),
    .D(_0821_),
    .Q(\dataMemory[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(net337),
    .D(_0822_),
    .Q(\dataMemory[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(net336),
    .D(_0823_),
    .Q(\dataMemory[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(net328),
    .D(_0824_),
    .Q(\dataMemory[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(net340),
    .D(_0825_),
    .Q(\dataMemory[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(net357),
    .D(_0826_),
    .Q(\dataMemory[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(net352),
    .D(_0827_),
    .Q(\dataMemory[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(net342),
    .D(_0828_),
    .Q(\dataMemory[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(net329),
    .D(_0829_),
    .Q(\dataMemory[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(net355),
    .D(_0830_),
    .Q(\dataMemory[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(net375),
    .D(_0831_),
    .Q(\dataMemory[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(net372),
    .D(_0832_),
    .Q(\dataMemory[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(net361),
    .D(_0833_),
    .Q(\dataMemory[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(net346),
    .D(_0834_),
    .Q(\dataMemory[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(net346),
    .D(_0835_),
    .Q(\dataMemory[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(net359),
    .D(_0836_),
    .Q(\dataMemory[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(net375),
    .D(_0837_),
    .Q(\dataMemory[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(net378),
    .D(_0838_),
    .Q(\dataMemory[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(net378),
    .D(_0839_),
    .Q(\dataMemory[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(net367),
    .D(_0840_),
    .Q(\dataMemory[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(net361),
    .D(_0841_),
    .Q(\dataMemory[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(net366),
    .D(_0842_),
    .Q(\dataMemory[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(net380),
    .D(_0843_),
    .Q(\dataMemory[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(net385),
    .D(_0844_),
    .Q(\dataMemory[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(net385),
    .D(_0845_),
    .Q(\dataMemory[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(net385),
    .D(_0846_),
    .Q(\dataMemory[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(net321),
    .D(_0847_),
    .Q(\dataMemory[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(net323),
    .D(_0848_),
    .Q(\dataMemory[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(net324),
    .D(_0849_),
    .Q(\dataMemory[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(net322),
    .D(_0850_),
    .Q(\dataMemory[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(net334),
    .D(_0851_),
    .Q(\dataMemory[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(net329),
    .D(_0852_),
    .Q(\dataMemory[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(net338),
    .D(_0853_),
    .Q(\dataMemory[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(net338),
    .D(_0854_),
    .Q(\dataMemory[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(net336),
    .D(_0855_),
    .Q(\dataMemory[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(net331),
    .D(_0856_),
    .Q(\dataMemory[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(net340),
    .D(_0857_),
    .Q(\dataMemory[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(net371),
    .D(_0858_),
    .Q(\dataMemory[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(net353),
    .D(_0859_),
    .Q(\dataMemory[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(net342),
    .D(_0860_),
    .Q(\dataMemory[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(net343),
    .D(_0861_),
    .Q(\dataMemory[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(net355),
    .D(_0862_),
    .Q(\dataMemory[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(net376),
    .D(_0863_),
    .Q(\dataMemory[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(net375),
    .D(_0864_),
    .Q(\dataMemory[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(net362),
    .D(_0865_),
    .Q(\dataMemory[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(net348),
    .D(_0866_),
    .Q(\dataMemory[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(net347),
    .D(_0867_),
    .Q(\dataMemory[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(net359),
    .D(_0868_),
    .Q(\dataMemory[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(net377),
    .D(_0869_),
    .Q(\dataMemory[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(net379),
    .D(_0870_),
    .Q(\dataMemory[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(net379),
    .D(_0871_),
    .Q(\dataMemory[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(net367),
    .D(_0872_),
    .Q(\dataMemory[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(net363),
    .D(_0873_),
    .Q(\dataMemory[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(net366),
    .D(_0874_),
    .Q(\dataMemory[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(net384),
    .D(_0875_),
    .Q(\dataMemory[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(net388),
    .D(_0876_),
    .Q(\dataMemory[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(net389),
    .D(_0877_),
    .Q(\dataMemory[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(net389),
    .D(_0878_),
    .Q(\dataMemory[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(net324),
    .D(_0879_),
    .Q(\dataMemory[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(net323),
    .D(_0880_),
    .Q(\dataMemory[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(net320),
    .D(_0881_),
    .Q(\dataMemory[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(net323),
    .D(_0882_),
    .Q(\dataMemory[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(net341),
    .D(_0883_),
    .Q(\dataMemory[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(net328),
    .D(_0884_),
    .Q(\dataMemory[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(net337),
    .D(_0885_),
    .Q(\dataMemory[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(net341),
    .D(_0886_),
    .Q(\dataMemory[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(net336),
    .D(_0887_),
    .Q(\dataMemory[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(net332),
    .D(_0888_),
    .Q(\dataMemory[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(net340),
    .D(_0889_),
    .Q(\dataMemory[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(net371),
    .D(_0890_),
    .Q(\dataMemory[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(net352),
    .D(_0891_),
    .Q(\dataMemory[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(net342),
    .D(_0892_),
    .Q(\dataMemory[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(net343),
    .D(_0893_),
    .Q(\dataMemory[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(net355),
    .D(_0894_),
    .Q(\dataMemory[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(net376),
    .D(_0895_),
    .Q(\dataMemory[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(net375),
    .D(_0896_),
    .Q(\dataMemory[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(net362),
    .D(_0897_),
    .Q(\dataMemory[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(net346),
    .D(_0898_),
    .Q(\dataMemory[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(net346),
    .D(_0899_),
    .Q(\dataMemory[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(net360),
    .D(_0900_),
    .Q(\dataMemory[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(net377),
    .D(_0901_),
    .Q(\dataMemory[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(net378),
    .D(_0902_),
    .Q(\dataMemory[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(net378),
    .D(_0903_),
    .Q(\dataMemory[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(net367),
    .D(_0904_),
    .Q(\dataMemory[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(net361),
    .D(_0905_),
    .Q(\dataMemory[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(net366),
    .D(_0906_),
    .Q(\dataMemory[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(net384),
    .D(_0907_),
    .Q(\dataMemory[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(net385),
    .D(_0908_),
    .Q(\dataMemory[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(net385),
    .D(_0909_),
    .Q(\dataMemory[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4632_ (.CLK(net385),
    .D(_0910_),
    .Q(\dataMemory[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(net316),
    .D(_0911_),
    .Q(\dataMemory[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(net323),
    .D(_0912_),
    .Q(\dataMemory[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(net320),
    .D(_0913_),
    .Q(\dataMemory[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(net323),
    .D(_0914_),
    .Q(\dataMemory[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(net341),
    .D(_0915_),
    .Q(\dataMemory[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(net328),
    .D(_0916_),
    .Q(\dataMemory[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(net334),
    .D(_0917_),
    .Q(\dataMemory[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(net337),
    .D(_0918_),
    .Q(\dataMemory[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(net336),
    .D(_0919_),
    .Q(\dataMemory[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(net328),
    .D(_0920_),
    .Q(\dataMemory[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4643_ (.CLK(net340),
    .D(_0921_),
    .Q(\dataMemory[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4644_ (.CLK(net360),
    .D(_0922_),
    .Q(\dataMemory[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(net341),
    .D(_0923_),
    .Q(\dataMemory[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(net343),
    .D(_0924_),
    .Q(\dataMemory[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4647_ (.CLK(net332),
    .D(_0925_),
    .Q(\dataMemory[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(net355),
    .D(_0926_),
    .Q(\dataMemory[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(net375),
    .D(_0927_),
    .Q(\dataMemory[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(net372),
    .D(_0928_),
    .Q(\dataMemory[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(net361),
    .D(_0929_),
    .Q(\dataMemory[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(net346),
    .D(_0930_),
    .Q(\dataMemory[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(net346),
    .D(_0931_),
    .Q(\dataMemory[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(net360),
    .D(_0932_),
    .Q(\dataMemory[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(net375),
    .D(_0933_),
    .Q(\dataMemory[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4656_ (.CLK(net378),
    .D(_0934_),
    .Q(\dataMemory[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4657_ (.CLK(net378),
    .D(_0935_),
    .Q(\dataMemory[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4658_ (.CLK(net366),
    .D(_0936_),
    .Q(\dataMemory[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(net347),
    .D(_0937_),
    .Q(\dataMemory[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4660_ (.CLK(net365),
    .D(_0938_),
    .Q(\dataMemory[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(net380),
    .D(_0939_),
    .Q(\dataMemory[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(net385),
    .D(_0940_),
    .Q(\dataMemory[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(net385),
    .D(_0941_),
    .Q(\dataMemory[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(net385),
    .D(_0942_),
    .Q(\dataMemory[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4665_ (.CLK(net320),
    .D(_0943_),
    .Q(\dataMemory[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4666_ (.CLK(net323),
    .D(_0944_),
    .Q(\dataMemory[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(net320),
    .D(_0945_),
    .Q(\dataMemory[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(net320),
    .D(_0946_),
    .Q(\dataMemory[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(net333),
    .D(_0947_),
    .Q(\dataMemory[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(net332),
    .D(_0948_),
    .Q(\dataMemory[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(net334),
    .D(_0949_),
    .Q(\dataMemory[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(net341),
    .D(_0950_),
    .Q(\dataMemory[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(net343),
    .D(_0951_),
    .Q(\dataMemory[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(net328),
    .D(_0952_),
    .Q(\dataMemory[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(net339),
    .D(_0953_),
    .Q(\dataMemory[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(net360),
    .D(_0954_),
    .Q(\dataMemory[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(net352),
    .D(_0955_),
    .Q(\dataMemory[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(net342),
    .D(_0956_),
    .Q(\dataMemory[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(net344),
    .D(_0957_),
    .Q(\dataMemory[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(net355),
    .D(_0958_),
    .Q(\dataMemory[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(net375),
    .D(_0959_),
    .Q(\dataMemory[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(net372),
    .D(_0960_),
    .Q(\dataMemory[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(net365),
    .D(_0961_),
    .Q(\dataMemory[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4684_ (.CLK(net350),
    .D(_0962_),
    .Q(\dataMemory[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(net350),
    .D(_0963_),
    .Q(\dataMemory[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(net360),
    .D(_0964_),
    .Q(\dataMemory[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(net377),
    .D(_0965_),
    .Q(\dataMemory[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(net378),
    .D(_0966_),
    .Q(\dataMemory[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4689_ (.CLK(net378),
    .D(_0967_),
    .Q(\dataMemory[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(net367),
    .D(_0968_),
    .Q(\dataMemory[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(net350),
    .D(_0969_),
    .Q(\dataMemory[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(net366),
    .D(_0970_),
    .Q(\dataMemory[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(net384),
    .D(_0971_),
    .Q(\dataMemory[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(net385),
    .D(_0972_),
    .Q(\dataMemory[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(net385),
    .D(_0973_),
    .Q(\dataMemory[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(net381),
    .D(_0974_),
    .Q(\dataMemory[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(net320),
    .D(_0975_),
    .Q(\dataMemory[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(net323),
    .D(_0976_),
    .Q(\dataMemory[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(net320),
    .D(_0977_),
    .Q(\dataMemory[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(net321),
    .D(_0978_),
    .Q(\dataMemory[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(net333),
    .D(_0979_),
    .Q(\dataMemory[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(net328),
    .D(_0980_),
    .Q(\dataMemory[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4703_ (.CLK(net334),
    .D(_0981_),
    .Q(\dataMemory[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(net337),
    .D(_0982_),
    .Q(\dataMemory[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(net343),
    .D(_0983_),
    .Q(\dataMemory[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(net329),
    .D(_0984_),
    .Q(\dataMemory[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(net339),
    .D(_0985_),
    .Q(\dataMemory[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(net360),
    .D(_0986_),
    .Q(\dataMemory[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(net352),
    .D(_0987_),
    .Q(\dataMemory[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(net345),
    .D(_0988_),
    .Q(\dataMemory[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(net344),
    .D(_0989_),
    .Q(\dataMemory[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(net354),
    .D(_0990_),
    .Q(\dataMemory[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(net375),
    .D(_0991_),
    .Q(\dataMemory[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(net372),
    .D(_0992_),
    .Q(\dataMemory[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(net362),
    .D(_0993_),
    .Q(\dataMemory[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(net345),
    .D(_0994_),
    .Q(\dataMemory[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(net348),
    .D(_0995_),
    .Q(\dataMemory[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(net358),
    .D(_0996_),
    .Q(\dataMemory[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(net377),
    .D(_0997_),
    .Q(\dataMemory[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4720_ (.CLK(net378),
    .D(_0998_),
    .Q(\dataMemory[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4721_ (.CLK(net378),
    .D(_0999_),
    .Q(\dataMemory[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4722_ (.CLK(net368),
    .D(_1000_),
    .Q(\dataMemory[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4723_ (.CLK(net350),
    .D(_1001_),
    .Q(\dataMemory[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4724_ (.CLK(net364),
    .D(_1002_),
    .Q(\dataMemory[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4725_ (.CLK(net384),
    .D(_1003_),
    .Q(\dataMemory[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4726_ (.CLK(net389),
    .D(_1004_),
    .Q(\dataMemory[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(net384),
    .D(_1005_),
    .Q(\dataMemory[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4728_ (.CLK(net381),
    .D(_1006_),
    .Q(\dataMemory[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4729_ (.CLK(net320),
    .D(_1007_),
    .Q(\dataMemory[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4730_ (.CLK(net323),
    .D(_1008_),
    .Q(\dataMemory[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4731_ (.CLK(net320),
    .D(_1009_),
    .Q(\dataMemory[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4732_ (.CLK(net321),
    .D(_1010_),
    .Q(\dataMemory[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4733_ (.CLK(net333),
    .D(_1011_),
    .Q(\dataMemory[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4734_ (.CLK(net328),
    .D(_1012_),
    .Q(\dataMemory[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4735_ (.CLK(net334),
    .D(_1013_),
    .Q(\dataMemory[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4736_ (.CLK(net337),
    .D(_1014_),
    .Q(\dataMemory[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4737_ (.CLK(net343),
    .D(_1015_),
    .Q(\dataMemory[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4738_ (.CLK(net329),
    .D(_1016_),
    .Q(\dataMemory[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4739_ (.CLK(net339),
    .D(_1017_),
    .Q(\dataMemory[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4740_ (.CLK(net360),
    .D(_1018_),
    .Q(\dataMemory[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4741_ (.CLK(net352),
    .D(_1019_),
    .Q(\dataMemory[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4742_ (.CLK(net343),
    .D(_1020_),
    .Q(\dataMemory[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4743_ (.CLK(net331),
    .D(_1021_),
    .Q(\dataMemory[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4744_ (.CLK(net354),
    .D(_1022_),
    .Q(\dataMemory[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4745_ (.CLK(net375),
    .D(_1023_),
    .Q(\dataMemory[14][16] ));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_16 fanout101 (.A(_1826_),
    .X(net101));
 sky130_fd_sc_hd__buf_8 fanout102 (.A(_1823_),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_1823_),
    .X(net103));
 sky130_fd_sc_hd__buf_8 fanout104 (.A(_1822_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_16 fanout105 (.A(_1822_),
    .X(net105));
 sky130_fd_sc_hd__buf_8 fanout106 (.A(_1821_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_16 fanout107 (.A(_1821_),
    .X(net107));
 sky130_fd_sc_hd__buf_8 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_16 fanout109 (.A(_1820_),
    .X(net109));
 sky130_fd_sc_hd__buf_8 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_12 fanout111 (.A(_1819_),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_16 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_16 fanout113 (.A(_1818_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_16 fanout115 (.A(_1817_),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_16 fanout117 (.A(_1815_),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout118 (.A(_1813_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_16 fanout119 (.A(_1813_),
    .X(net119));
 sky130_fd_sc_hd__buf_8 fanout120 (.A(_1812_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_16 fanout121 (.A(_1812_),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(_1809_),
    .X(net122));
 sky130_fd_sc_hd__buf_8 fanout123 (.A(_1809_),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_16 fanout125 (.A(_1802_),
    .X(net125));
 sky130_fd_sc_hd__buf_8 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_16 fanout127 (.A(_1843_),
    .X(net127));
 sky130_fd_sc_hd__buf_8 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_16 fanout129 (.A(_1838_),
    .X(net129));
 sky130_fd_sc_hd__buf_8 fanout130 (.A(_1835_),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_16 fanout131 (.A(_1835_),
    .X(net131));
 sky130_fd_sc_hd__buf_8 fanout132 (.A(_1824_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_16 fanout133 (.A(_1824_),
    .X(net133));
 sky130_fd_sc_hd__buf_8 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_16 fanout135 (.A(_1805_),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net150),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net150),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net150),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net150),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 fanout140 (.A(net142),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_8 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_8 fanout142 (.A(net150),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net145),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_6 fanout145 (.A(net150),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_8 fanout146 (.A(net150),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 fanout147 (.A(net150),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_8 fanout148 (.A(net150),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_8 fanout150 (.A(_1028_),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_8 fanout151 (.A(net166),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net166),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_8 fanout153 (.A(net166),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(net166),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_8 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(net166),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_8 fanout158 (.A(net161),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_8 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net166),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net166),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(net166),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net166),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(_1027_),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_8 fanout167 (.A(net182),
    .X(net167));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net182),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net182),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(net182),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_8 fanout171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_8 fanout173 (.A(net182),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 fanout174 (.A(net177),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net177),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(net182),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_4 fanout179 (.A(net182),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_6 fanout182 (.A(_1026_),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(_1025_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_8 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_8 fanout186 (.A(_1025_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_8 fanout187 (.A(net196),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net196),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(net196),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(net196),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net195),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_8 fanout192 (.A(net195),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_8 fanout193 (.A(net195),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_8 fanout196 (.A(_1024_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 fanout197 (.A(net9),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(net9),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 fanout200 (.A(net8),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net7),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_16 fanout203 (.A(net205),
    .X(net203));
 sky130_fd_sc_hd__buf_8 fanout204 (.A(net205),
    .X(net204));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(net6),
    .X(net205));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_8 fanout207 (.A(net210),
    .X(net207));
 sky130_fd_sc_hd__buf_6 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_6 fanout210 (.A(net5),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net215),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net215),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_8 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net221),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_8 fanout216 (.A(net221),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(net221),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net221),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_8 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_6 fanout221 (.A(net4),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(net38),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net37),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_4 fanout225 (.A(net37),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net36),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(net35),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net35),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net34),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net33),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net32),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 fanout235 (.A(net32),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net31),
    .X(net236));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(net31),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_4 fanout239 (.A(net30),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net248),
    .X(net240));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net248),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net248),
    .X(net242));
 sky130_fd_sc_hd__buf_4 fanout243 (.A(net248),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(net248),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(net3),
    .X(net248));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(net3),
    .X(net249));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net3),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net3),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(net257),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net257),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(net3),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net29),
    .X(net259));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(net28),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 fanout262 (.A(net27),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 fanout263 (.A(net27),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(net26),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net26),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_4 fanout267 (.A(net25),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net24),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net23),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(net22),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net21),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net21),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net20),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(net20),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_8 fanout279 (.A(net286),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net286),
    .X(net280));
 sky130_fd_sc_hd__buf_4 fanout281 (.A(net286),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_8 fanout283 (.A(net286),
    .X(net283));
 sky130_fd_sc_hd__buf_4 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_8 fanout286 (.A(net2),
    .X(net286));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_8 fanout288 (.A(net2),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(net2),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net2),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 fanout291 (.A(net295),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(net295),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_8 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(net2),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net19),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 fanout297 (.A(net19),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 fanout298 (.A(net18),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(net18),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_4 fanout301 (.A(net17),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(net16),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_4 fanout303 (.A(net16),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net15),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(net15),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 fanout306 (.A(net14),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(net14),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 fanout309 (.A(net13),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_4 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 fanout311 (.A(net12),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 fanout312 (.A(net11),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(net11),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net10),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(net10),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_4 fanout317 (.A(net324),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 fanout318 (.A(net324),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 fanout319 (.A(net324),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(net324),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 fanout324 (.A(net332),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 fanout327 (.A(net332),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_4 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_4 fanout329 (.A(net332),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_4 fanout330 (.A(net332),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 fanout331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 fanout332 (.A(net351),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 fanout333 (.A(net341),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 fanout334 (.A(net341),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_4 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_4 fanout336 (.A(net341),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(net341),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 fanout339 (.A(net341),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(net351),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 fanout343 (.A(net351),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_4 fanout344 (.A(net351),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 fanout345 (.A(net351),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 fanout346 (.A(net350),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 fanout347 (.A(net350),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_4 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__buf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_4 fanout351 (.A(net1),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_4 fanout353 (.A(net370),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 fanout354 (.A(net370),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_4 fanout355 (.A(net370),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 fanout356 (.A(net357),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 fanout357 (.A(net360),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_4 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_4 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_2 fanout360 (.A(net370),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_4 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__buf_4 fanout362 (.A(net365),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 fanout363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_2 fanout365 (.A(net370),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_4 fanout366 (.A(net370),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(net370),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_4 fanout370 (.A(net1),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(net390),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_4 fanout372 (.A(net390),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_4 fanout373 (.A(net390),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_4 fanout374 (.A(net390),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net377),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(net390),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_4 fanout378 (.A(net390),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_4 fanout379 (.A(net390),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_4 fanout380 (.A(net384),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_4 fanout381 (.A(net384),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(net384),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_4 fanout384 (.A(net389),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_4 fanout385 (.A(net389),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_4 fanout386 (.A(net389),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_4 fanout387 (.A(net389),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_4 fanout388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_4 fanout390 (.A(net1),
    .X(net390));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_16 fanout73 (.A(_1844_),
    .X(net73));
 sky130_fd_sc_hd__buf_8 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(_1842_),
    .X(net75));
 sky130_fd_sc_hd__buf_8 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_16 fanout77 (.A(_1841_),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(_1840_),
    .X(net79));
 sky130_fd_sc_hd__buf_8 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_8 fanout81 (.A(_1839_),
    .X(net81));
 sky130_fd_sc_hd__buf_8 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_16 fanout83 (.A(_1837_),
    .X(net83));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_16 fanout85 (.A(_1836_),
    .X(net85));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_16 fanout87 (.A(_1834_),
    .X(net87));
 sky130_fd_sc_hd__buf_8 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_16 fanout89 (.A(_1833_),
    .X(net89));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_16 fanout91 (.A(_1832_),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_12 fanout93 (.A(_1831_),
    .X(net93));
 sky130_fd_sc_hd__buf_8 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(_1830_),
    .X(net95));
 sky130_fd_sc_hd__buf_8 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_16 fanout97 (.A(_1828_),
    .X(net97));
 sky130_fd_sc_hd__buf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_12 fanout99 (.A(_1827_),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(clock),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(dataMemDataP2M[12]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(dataMemDataP2M[13]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(dataMemDataP2M[14]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(dataMemDataP2M[15]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(dataMemDataP2M[16]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(dataMemDataP2M[17]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(dataMemDataP2M[18]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(dataMemDataP2M[19]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(dataMemDataP2M[1]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(dataMemDataP2M[20]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(dataMemAddr[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(dataMemDataP2M[21]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(dataMemDataP2M[22]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(dataMemDataP2M[23]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(dataMemDataP2M[24]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(dataMemDataP2M[25]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(dataMemDataP2M[26]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(dataMemDataP2M[27]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(dataMemDataP2M[28]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(dataMemDataP2M[29]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(dataMemDataP2M[2]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(dataMemAddr[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(dataMemDataP2M[30]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(dataMemDataP2M[31]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(dataMemDataP2M[3]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(dataMemDataP2M[4]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(dataMemDataP2M[5]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(dataMemDataP2M[6]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(dataMemDataP2M[7]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(dataMemDataP2M[8]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(dataMemDataP2M[9]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(dataMemWen),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(dataMemAddr[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(dataMemAddr[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(dataMemAddr[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(dataMemDataP2M[0]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(dataMemDataP2M[10]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(dataMemDataP2M[11]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(dataMemDataM2P[0]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(dataMemDataM2P[10]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(dataMemDataM2P[11]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(dataMemDataM2P[12]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(dataMemDataM2P[13]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(dataMemDataM2P[14]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(dataMemDataM2P[15]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(dataMemDataM2P[16]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(dataMemDataM2P[17]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(dataMemDataM2P[18]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(dataMemDataM2P[19]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(dataMemDataM2P[1]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(dataMemDataM2P[20]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(dataMemDataM2P[21]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(dataMemDataM2P[22]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(dataMemDataM2P[23]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(dataMemDataM2P[24]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(dataMemDataM2P[25]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(dataMemDataM2P[26]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(dataMemDataM2P[27]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(dataMemDataM2P[28]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net61),
    .X(dataMemDataM2P[29]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(dataMemDataM2P[2]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(dataMemDataM2P[30]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(dataMemDataM2P[31]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(dataMemDataM2P[3]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(dataMemDataM2P[4]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(dataMemDataM2P[5]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(dataMemDataM2P[6]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(dataMemDataM2P[7]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(dataMemDataM2P[8]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(dataMemDataM2P[9]));
endmodule

